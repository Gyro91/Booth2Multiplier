

library IEEE;
use IEEE.std_logic_1164.all;

entity booth2_tbn8 IS

end booth2_tbn8;

-- Test Booth multiplier for N=M=8

architecture booth2_tbn8 of booth2_tbn8 is
	component Booth2Multiplier
  	generic(N : integer := 4; 
            M : integer := 4   
       );
	port (
	x : in  std_logic_vector(N-1 downto 0); 	-- x is the multiplicand
	y : in  std_logic_vector(M-1 downto 0);		-- y is the multiplier
	z : out	std_logic_vector(N+M-1 downto 0)	-- z is the result of the multiplication
		);
	end component; 
	
   constant MckPer  :  time     := 200 ns;  -- Master Clk period
	   
   signal   clk  : std_logic := '0';
   signal   x_in   	: std_logic_VECTOR (7 downto 0):="00000000";
   signal   y_in    : std_logic_VECTOR (7 downto 0):="00000000";	
   signal   z_out   : std_logic_VECTOR (15 downto 0):="0000000000000000";
   signal clk_cycle : integer;
   signal Testing: boolean := True;	
   signal  z_correct   : std_logic_VECTOR (15 downto 0):="0000000000000000";
   signal 	diff		: std_logic := '0';
begin 			 
	I: Booth2Multiplier generic map(N=>8, M=>8)
		port map(x=>x_in,y=>y_in, z=>z_out);
				
		clk <= not clk after MckPer/2 when Testing else '0';


   Test_Proc: process(clk)
   variable count: INTEGER:= 0;
   
   begin
     clk_cycle <= (count+1)/2;

     case clk_cycle is
                  when 0 => y_in <= "10000000"; x_in <= "10000000"; z_correct<="0100000000000000";
        when 1 => y_in <= "10000000"; x_in <= "10000001"; z_correct<="0011111110000000";
        when 2 => y_in <= "10000000"; x_in <= "10000010"; z_correct<="0011111100000000";
        when 3 => y_in <= "10000000"; x_in <= "10000011"; z_correct<="0011111010000000";
        when 4 => y_in <= "10000000"; x_in <= "10000100"; z_correct<="0011111000000000";
        when 5 => y_in <= "10000000"; x_in <= "10000101"; z_correct<="0011110110000000";
        when 6 => y_in <= "10000000"; x_in <= "10000110"; z_correct<="0011110100000000";
        when 7 => y_in <= "10000000"; x_in <= "10000111"; z_correct<="0011110010000000";
        when 8 => y_in <= "10000000"; x_in <= "10001000"; z_correct<="0011110000000000";
        when 9 => y_in <= "10000000"; x_in <= "10001001"; z_correct<="0011101110000000";
        when 10 => y_in <= "10000000"; x_in <= "10001010"; z_correct<="0011101100000000";
        when 11 => y_in <= "10000000"; x_in <= "10001011"; z_correct<="0011101010000000";
        when 12 => y_in <= "10000000"; x_in <= "10001100"; z_correct<="0011101000000000";
        when 13 => y_in <= "10000000"; x_in <= "10001101"; z_correct<="0011100110000000";
        when 14 => y_in <= "10000000"; x_in <= "10001110"; z_correct<="0011100100000000";
        when 15 => y_in <= "10000000"; x_in <= "10001111"; z_correct<="0011100010000000";
        when 16 => y_in <= "10000000"; x_in <= "10010000"; z_correct<="0011100000000000";
        when 17 => y_in <= "10000000"; x_in <= "10010001"; z_correct<="0011011110000000";
        when 18 => y_in <= "10000000"; x_in <= "10010010"; z_correct<="0011011100000000";
        when 19 => y_in <= "10000000"; x_in <= "10010011"; z_correct<="0011011010000000";
        when 20 => y_in <= "10000000"; x_in <= "10010100"; z_correct<="0011011000000000";
        when 21 => y_in <= "10000000"; x_in <= "10010101"; z_correct<="0011010110000000";
        when 22 => y_in <= "10000000"; x_in <= "10010110"; z_correct<="0011010100000000";
        when 23 => y_in <= "10000000"; x_in <= "10010111"; z_correct<="0011010010000000";
        when 24 => y_in <= "10000000"; x_in <= "10011000"; z_correct<="0011010000000000";
        when 25 => y_in <= "10000000"; x_in <= "10011001"; z_correct<="0011001110000000";
        when 26 => y_in <= "10000000"; x_in <= "10011010"; z_correct<="0011001100000000";
        when 27 => y_in <= "10000000"; x_in <= "10011011"; z_correct<="0011001010000000";
        when 28 => y_in <= "10000000"; x_in <= "10011100"; z_correct<="0011001000000000";
        when 29 => y_in <= "10000000"; x_in <= "10011101"; z_correct<="0011000110000000";
        when 30 => y_in <= "10000000"; x_in <= "10011110"; z_correct<="0011000100000000";
        when 31 => y_in <= "10000000"; x_in <= "10011111"; z_correct<="0011000010000000";
        when 32 => y_in <= "10000000"; x_in <= "10100000"; z_correct<="0011000000000000";
        when 33 => y_in <= "10000000"; x_in <= "10100001"; z_correct<="0010111110000000";
        when 34 => y_in <= "10000000"; x_in <= "10100010"; z_correct<="0010111100000000";
        when 35 => y_in <= "10000000"; x_in <= "10100011"; z_correct<="0010111010000000";
        when 36 => y_in <= "10000000"; x_in <= "10100100"; z_correct<="0010111000000000";
        when 37 => y_in <= "10000000"; x_in <= "10100101"; z_correct<="0010110110000000";
        when 38 => y_in <= "10000000"; x_in <= "10100110"; z_correct<="0010110100000000";
        when 39 => y_in <= "10000000"; x_in <= "10100111"; z_correct<="0010110010000000";
        when 40 => y_in <= "10000000"; x_in <= "10101000"; z_correct<="0010110000000000";
        when 41 => y_in <= "10000000"; x_in <= "10101001"; z_correct<="0010101110000000";
        when 42 => y_in <= "10000000"; x_in <= "10101010"; z_correct<="0010101100000000";
        when 43 => y_in <= "10000000"; x_in <= "10101011"; z_correct<="0010101010000000";
        when 44 => y_in <= "10000000"; x_in <= "10101100"; z_correct<="0010101000000000";
        when 45 => y_in <= "10000000"; x_in <= "10101101"; z_correct<="0010100110000000";
        when 46 => y_in <= "10000000"; x_in <= "10101110"; z_correct<="0010100100000000";
        when 47 => y_in <= "10000000"; x_in <= "10101111"; z_correct<="0010100010000000";
        when 48 => y_in <= "10000000"; x_in <= "10110000"; z_correct<="0010100000000000";
        when 49 => y_in <= "10000000"; x_in <= "10110001"; z_correct<="0010011110000000";
        when 50 => y_in <= "10000000"; x_in <= "10110010"; z_correct<="0010011100000000";
        when 51 => y_in <= "10000000"; x_in <= "10110011"; z_correct<="0010011010000000";
        when 52 => y_in <= "10000000"; x_in <= "10110100"; z_correct<="0010011000000000";
        when 53 => y_in <= "10000000"; x_in <= "10110101"; z_correct<="0010010110000000";
        when 54 => y_in <= "10000000"; x_in <= "10110110"; z_correct<="0010010100000000";
        when 55 => y_in <= "10000000"; x_in <= "10110111"; z_correct<="0010010010000000";
        when 56 => y_in <= "10000000"; x_in <= "10111000"; z_correct<="0010010000000000";
        when 57 => y_in <= "10000000"; x_in <= "10111001"; z_correct<="0010001110000000";
        when 58 => y_in <= "10000000"; x_in <= "10111010"; z_correct<="0010001100000000";
        when 59 => y_in <= "10000000"; x_in <= "10111011"; z_correct<="0010001010000000";
        when 60 => y_in <= "10000000"; x_in <= "10111100"; z_correct<="0010001000000000";
        when 61 => y_in <= "10000000"; x_in <= "10111101"; z_correct<="0010000110000000";
        when 62 => y_in <= "10000000"; x_in <= "10111110"; z_correct<="0010000100000000";
        when 63 => y_in <= "10000000"; x_in <= "10111111"; z_correct<="0010000010000000";
        when 64 => y_in <= "10000000"; x_in <= "11000000"; z_correct<="0010000000000000";
        when 65 => y_in <= "10000000"; x_in <= "11000001"; z_correct<="0001111110000000";
        when 66 => y_in <= "10000000"; x_in <= "11000010"; z_correct<="0001111100000000";
        when 67 => y_in <= "10000000"; x_in <= "11000011"; z_correct<="0001111010000000";
        when 68 => y_in <= "10000000"; x_in <= "11000100"; z_correct<="0001111000000000";
        when 69 => y_in <= "10000000"; x_in <= "11000101"; z_correct<="0001110110000000";
        when 70 => y_in <= "10000000"; x_in <= "11000110"; z_correct<="0001110100000000";
        when 71 => y_in <= "10000000"; x_in <= "11000111"; z_correct<="0001110010000000";
        when 72 => y_in <= "10000000"; x_in <= "11001000"; z_correct<="0001110000000000";
        when 73 => y_in <= "10000000"; x_in <= "11001001"; z_correct<="0001101110000000";
        when 74 => y_in <= "10000000"; x_in <= "11001010"; z_correct<="0001101100000000";
        when 75 => y_in <= "10000000"; x_in <= "11001011"; z_correct<="0001101010000000";
        when 76 => y_in <= "10000000"; x_in <= "11001100"; z_correct<="0001101000000000";
        when 77 => y_in <= "10000000"; x_in <= "11001101"; z_correct<="0001100110000000";
        when 78 => y_in <= "10000000"; x_in <= "11001110"; z_correct<="0001100100000000";
        when 79 => y_in <= "10000000"; x_in <= "11001111"; z_correct<="0001100010000000";
        when 80 => y_in <= "10000000"; x_in <= "11010000"; z_correct<="0001100000000000";
        when 81 => y_in <= "10000000"; x_in <= "11010001"; z_correct<="0001011110000000";
        when 82 => y_in <= "10000000"; x_in <= "11010010"; z_correct<="0001011100000000";
        when 83 => y_in <= "10000000"; x_in <= "11010011"; z_correct<="0001011010000000";
        when 84 => y_in <= "10000000"; x_in <= "11010100"; z_correct<="0001011000000000";
        when 85 => y_in <= "10000000"; x_in <= "11010101"; z_correct<="0001010110000000";
        when 86 => y_in <= "10000000"; x_in <= "11010110"; z_correct<="0001010100000000";
        when 87 => y_in <= "10000000"; x_in <= "11010111"; z_correct<="0001010010000000";
        when 88 => y_in <= "10000000"; x_in <= "11011000"; z_correct<="0001010000000000";
        when 89 => y_in <= "10000000"; x_in <= "11011001"; z_correct<="0001001110000000";
        when 90 => y_in <= "10000000"; x_in <= "11011010"; z_correct<="0001001100000000";
        when 91 => y_in <= "10000000"; x_in <= "11011011"; z_correct<="0001001010000000";
        when 92 => y_in <= "10000000"; x_in <= "11011100"; z_correct<="0001001000000000";
        when 93 => y_in <= "10000000"; x_in <= "11011101"; z_correct<="0001000110000000";
        when 94 => y_in <= "10000000"; x_in <= "11011110"; z_correct<="0001000100000000";
        when 95 => y_in <= "10000000"; x_in <= "11011111"; z_correct<="0001000010000000";
        when 96 => y_in <= "10000000"; x_in <= "11100000"; z_correct<="0001000000000000";
        when 97 => y_in <= "10000000"; x_in <= "11100001"; z_correct<="0000111110000000";
        when 98 => y_in <= "10000000"; x_in <= "11100010"; z_correct<="0000111100000000";
        when 99 => y_in <= "10000000"; x_in <= "11100011"; z_correct<="0000111010000000";
        when 100 => y_in <= "10000000"; x_in <= "11100100"; z_correct<="0000111000000000";
        when 101 => y_in <= "10000000"; x_in <= "11100101"; z_correct<="0000110110000000";
        when 102 => y_in <= "10000000"; x_in <= "11100110"; z_correct<="0000110100000000";
        when 103 => y_in <= "10000000"; x_in <= "11100111"; z_correct<="0000110010000000";
        when 104 => y_in <= "10000000"; x_in <= "11101000"; z_correct<="0000110000000000";
        when 105 => y_in <= "10000000"; x_in <= "11101001"; z_correct<="0000101110000000";
        when 106 => y_in <= "10000000"; x_in <= "11101010"; z_correct<="0000101100000000";
        when 107 => y_in <= "10000000"; x_in <= "11101011"; z_correct<="0000101010000000";
        when 108 => y_in <= "10000000"; x_in <= "11101100"; z_correct<="0000101000000000";
        when 109 => y_in <= "10000000"; x_in <= "11101101"; z_correct<="0000100110000000";
        when 110 => y_in <= "10000000"; x_in <= "11101110"; z_correct<="0000100100000000";
        when 111 => y_in <= "10000000"; x_in <= "11101111"; z_correct<="0000100010000000";
        when 112 => y_in <= "10000000"; x_in <= "11110000"; z_correct<="0000100000000000";
        when 113 => y_in <= "10000000"; x_in <= "11110001"; z_correct<="0000011110000000";
        when 114 => y_in <= "10000000"; x_in <= "11110010"; z_correct<="0000011100000000";
        when 115 => y_in <= "10000000"; x_in <= "11110011"; z_correct<="0000011010000000";
        when 116 => y_in <= "10000000"; x_in <= "11110100"; z_correct<="0000011000000000";
        when 117 => y_in <= "10000000"; x_in <= "11110101"; z_correct<="0000010110000000";
        when 118 => y_in <= "10000000"; x_in <= "11110110"; z_correct<="0000010100000000";
        when 119 => y_in <= "10000000"; x_in <= "11110111"; z_correct<="0000010010000000";
        when 120 => y_in <= "10000000"; x_in <= "11111000"; z_correct<="0000010000000000";
        when 121 => y_in <= "10000000"; x_in <= "11111001"; z_correct<="0000001110000000";
        when 122 => y_in <= "10000000"; x_in <= "11111010"; z_correct<="0000001100000000";
        when 123 => y_in <= "10000000"; x_in <= "11111011"; z_correct<="0000001010000000";
        when 124 => y_in <= "10000000"; x_in <= "11111100"; z_correct<="0000001000000000";
        when 125 => y_in <= "10000000"; x_in <= "11111101"; z_correct<="0000000110000000";
        when 126 => y_in <= "10000000"; x_in <= "11111110"; z_correct<="0000000100000000";
        when 127 => y_in <= "10000000"; x_in <= "11111111"; z_correct<="0000000010000000";
        when 128 => y_in <= "10000000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 129 => y_in <= "10000000"; x_in <= "00000001"; z_correct<="1111111110000000";
        when 130 => y_in <= "10000000"; x_in <= "00000010"; z_correct<="1111111100000000";
        when 131 => y_in <= "10000000"; x_in <= "00000011"; z_correct<="1111111010000000";
        when 132 => y_in <= "10000000"; x_in <= "00000100"; z_correct<="1111111000000000";
        when 133 => y_in <= "10000000"; x_in <= "00000101"; z_correct<="1111110110000000";
        when 134 => y_in <= "10000000"; x_in <= "00000110"; z_correct<="1111110100000000";
        when 135 => y_in <= "10000000"; x_in <= "00000111"; z_correct<="1111110010000000";
        when 136 => y_in <= "10000000"; x_in <= "00001000"; z_correct<="1111110000000000";
        when 137 => y_in <= "10000000"; x_in <= "00001001"; z_correct<="1111101110000000";
        when 138 => y_in <= "10000000"; x_in <= "00001010"; z_correct<="1111101100000000";
        when 139 => y_in <= "10000000"; x_in <= "00001011"; z_correct<="1111101010000000";
        when 140 => y_in <= "10000000"; x_in <= "00001100"; z_correct<="1111101000000000";
        when 141 => y_in <= "10000000"; x_in <= "00001101"; z_correct<="1111100110000000";
        when 142 => y_in <= "10000000"; x_in <= "00001110"; z_correct<="1111100100000000";
        when 143 => y_in <= "10000000"; x_in <= "00001111"; z_correct<="1111100010000000";
        when 144 => y_in <= "10000000"; x_in <= "00010000"; z_correct<="1111100000000000";
        when 145 => y_in <= "10000000"; x_in <= "00010001"; z_correct<="1111011110000000";
        when 146 => y_in <= "10000000"; x_in <= "00010010"; z_correct<="1111011100000000";
        when 147 => y_in <= "10000000"; x_in <= "00010011"; z_correct<="1111011010000000";
        when 148 => y_in <= "10000000"; x_in <= "00010100"; z_correct<="1111011000000000";
        when 149 => y_in <= "10000000"; x_in <= "00010101"; z_correct<="1111010110000000";
        when 150 => y_in <= "10000000"; x_in <= "00010110"; z_correct<="1111010100000000";
        when 151 => y_in <= "10000000"; x_in <= "00010111"; z_correct<="1111010010000000";
        when 152 => y_in <= "10000000"; x_in <= "00011000"; z_correct<="1111010000000000";
        when 153 => y_in <= "10000000"; x_in <= "00011001"; z_correct<="1111001110000000";
        when 154 => y_in <= "10000000"; x_in <= "00011010"; z_correct<="1111001100000000";
        when 155 => y_in <= "10000000"; x_in <= "00011011"; z_correct<="1111001010000000";
        when 156 => y_in <= "10000000"; x_in <= "00011100"; z_correct<="1111001000000000";
        when 157 => y_in <= "10000000"; x_in <= "00011101"; z_correct<="1111000110000000";
        when 158 => y_in <= "10000000"; x_in <= "00011110"; z_correct<="1111000100000000";
        when 159 => y_in <= "10000000"; x_in <= "00011111"; z_correct<="1111000010000000";
        when 160 => y_in <= "10000000"; x_in <= "00100000"; z_correct<="1111000000000000";
        when 161 => y_in <= "10000000"; x_in <= "00100001"; z_correct<="1110111110000000";
        when 162 => y_in <= "10000000"; x_in <= "00100010"; z_correct<="1110111100000000";
        when 163 => y_in <= "10000000"; x_in <= "00100011"; z_correct<="1110111010000000";
        when 164 => y_in <= "10000000"; x_in <= "00100100"; z_correct<="1110111000000000";
        when 165 => y_in <= "10000000"; x_in <= "00100101"; z_correct<="1110110110000000";
        when 166 => y_in <= "10000000"; x_in <= "00100110"; z_correct<="1110110100000000";
        when 167 => y_in <= "10000000"; x_in <= "00100111"; z_correct<="1110110010000000";
        when 168 => y_in <= "10000000"; x_in <= "00101000"; z_correct<="1110110000000000";
        when 169 => y_in <= "10000000"; x_in <= "00101001"; z_correct<="1110101110000000";
        when 170 => y_in <= "10000000"; x_in <= "00101010"; z_correct<="1110101100000000";
        when 171 => y_in <= "10000000"; x_in <= "00101011"; z_correct<="1110101010000000";
        when 172 => y_in <= "10000000"; x_in <= "00101100"; z_correct<="1110101000000000";
        when 173 => y_in <= "10000000"; x_in <= "00101101"; z_correct<="1110100110000000";
        when 174 => y_in <= "10000000"; x_in <= "00101110"; z_correct<="1110100100000000";
        when 175 => y_in <= "10000000"; x_in <= "00101111"; z_correct<="1110100010000000";
        when 176 => y_in <= "10000000"; x_in <= "00110000"; z_correct<="1110100000000000";
        when 177 => y_in <= "10000000"; x_in <= "00110001"; z_correct<="1110011110000000";
        when 178 => y_in <= "10000000"; x_in <= "00110010"; z_correct<="1110011100000000";
        when 179 => y_in <= "10000000"; x_in <= "00110011"; z_correct<="1110011010000000";
        when 180 => y_in <= "10000000"; x_in <= "00110100"; z_correct<="1110011000000000";
        when 181 => y_in <= "10000000"; x_in <= "00110101"; z_correct<="1110010110000000";
        when 182 => y_in <= "10000000"; x_in <= "00110110"; z_correct<="1110010100000000";
        when 183 => y_in <= "10000000"; x_in <= "00110111"; z_correct<="1110010010000000";
        when 184 => y_in <= "10000000"; x_in <= "00111000"; z_correct<="1110010000000000";
        when 185 => y_in <= "10000000"; x_in <= "00111001"; z_correct<="1110001110000000";
        when 186 => y_in <= "10000000"; x_in <= "00111010"; z_correct<="1110001100000000";
        when 187 => y_in <= "10000000"; x_in <= "00111011"; z_correct<="1110001010000000";
        when 188 => y_in <= "10000000"; x_in <= "00111100"; z_correct<="1110001000000000";
        when 189 => y_in <= "10000000"; x_in <= "00111101"; z_correct<="1110000110000000";
        when 190 => y_in <= "10000000"; x_in <= "00111110"; z_correct<="1110000100000000";
        when 191 => y_in <= "10000000"; x_in <= "00111111"; z_correct<="1110000010000000";
        when 192 => y_in <= "10000000"; x_in <= "01000000"; z_correct<="1110000000000000";
        when 193 => y_in <= "10000000"; x_in <= "01000001"; z_correct<="1101111110000000";
        when 194 => y_in <= "10000000"; x_in <= "01000010"; z_correct<="1101111100000000";
        when 195 => y_in <= "10000000"; x_in <= "01000011"; z_correct<="1101111010000000";
        when 196 => y_in <= "10000000"; x_in <= "01000100"; z_correct<="1101111000000000";
        when 197 => y_in <= "10000000"; x_in <= "01000101"; z_correct<="1101110110000000";
        when 198 => y_in <= "10000000"; x_in <= "01000110"; z_correct<="1101110100000000";
        when 199 => y_in <= "10000000"; x_in <= "01000111"; z_correct<="1101110010000000";
        when 200 => y_in <= "10000000"; x_in <= "01001000"; z_correct<="1101110000000000";
        when 201 => y_in <= "10000000"; x_in <= "01001001"; z_correct<="1101101110000000";
        when 202 => y_in <= "10000000"; x_in <= "01001010"; z_correct<="1101101100000000";
        when 203 => y_in <= "10000000"; x_in <= "01001011"; z_correct<="1101101010000000";
        when 204 => y_in <= "10000000"; x_in <= "01001100"; z_correct<="1101101000000000";
        when 205 => y_in <= "10000000"; x_in <= "01001101"; z_correct<="1101100110000000";
        when 206 => y_in <= "10000000"; x_in <= "01001110"; z_correct<="1101100100000000";
        when 207 => y_in <= "10000000"; x_in <= "01001111"; z_correct<="1101100010000000";
        when 208 => y_in <= "10000000"; x_in <= "01010000"; z_correct<="1101100000000000";
        when 209 => y_in <= "10000000"; x_in <= "01010001"; z_correct<="1101011110000000";
        when 210 => y_in <= "10000000"; x_in <= "01010010"; z_correct<="1101011100000000";
        when 211 => y_in <= "10000000"; x_in <= "01010011"; z_correct<="1101011010000000";
        when 212 => y_in <= "10000000"; x_in <= "01010100"; z_correct<="1101011000000000";
        when 213 => y_in <= "10000000"; x_in <= "01010101"; z_correct<="1101010110000000";
        when 214 => y_in <= "10000000"; x_in <= "01010110"; z_correct<="1101010100000000";
        when 215 => y_in <= "10000000"; x_in <= "01010111"; z_correct<="1101010010000000";
        when 216 => y_in <= "10000000"; x_in <= "01011000"; z_correct<="1101010000000000";
        when 217 => y_in <= "10000000"; x_in <= "01011001"; z_correct<="1101001110000000";
        when 218 => y_in <= "10000000"; x_in <= "01011010"; z_correct<="1101001100000000";
        when 219 => y_in <= "10000000"; x_in <= "01011011"; z_correct<="1101001010000000";
        when 220 => y_in <= "10000000"; x_in <= "01011100"; z_correct<="1101001000000000";
        when 221 => y_in <= "10000000"; x_in <= "01011101"; z_correct<="1101000110000000";
        when 222 => y_in <= "10000000"; x_in <= "01011110"; z_correct<="1101000100000000";
        when 223 => y_in <= "10000000"; x_in <= "01011111"; z_correct<="1101000010000000";
        when 224 => y_in <= "10000000"; x_in <= "01100000"; z_correct<="1101000000000000";
        when 225 => y_in <= "10000000"; x_in <= "01100001"; z_correct<="1100111110000000";
        when 226 => y_in <= "10000000"; x_in <= "01100010"; z_correct<="1100111100000000";
        when 227 => y_in <= "10000000"; x_in <= "01100011"; z_correct<="1100111010000000";
        when 228 => y_in <= "10000000"; x_in <= "01100100"; z_correct<="1100111000000000";
        when 229 => y_in <= "10000000"; x_in <= "01100101"; z_correct<="1100110110000000";
        when 230 => y_in <= "10000000"; x_in <= "01100110"; z_correct<="1100110100000000";
        when 231 => y_in <= "10000000"; x_in <= "01100111"; z_correct<="1100110010000000";
        when 232 => y_in <= "10000000"; x_in <= "01101000"; z_correct<="1100110000000000";
        when 233 => y_in <= "10000000"; x_in <= "01101001"; z_correct<="1100101110000000";
        when 234 => y_in <= "10000000"; x_in <= "01101010"; z_correct<="1100101100000000";
        when 235 => y_in <= "10000000"; x_in <= "01101011"; z_correct<="1100101010000000";
        when 236 => y_in <= "10000000"; x_in <= "01101100"; z_correct<="1100101000000000";
        when 237 => y_in <= "10000000"; x_in <= "01101101"; z_correct<="1100100110000000";
        when 238 => y_in <= "10000000"; x_in <= "01101110"; z_correct<="1100100100000000";
        when 239 => y_in <= "10000000"; x_in <= "01101111"; z_correct<="1100100010000000";
        when 240 => y_in <= "10000000"; x_in <= "01110000"; z_correct<="1100100000000000";
        when 241 => y_in <= "10000000"; x_in <= "01110001"; z_correct<="1100011110000000";
        when 242 => y_in <= "10000000"; x_in <= "01110010"; z_correct<="1100011100000000";
        when 243 => y_in <= "10000000"; x_in <= "01110011"; z_correct<="1100011010000000";
        when 244 => y_in <= "10000000"; x_in <= "01110100"; z_correct<="1100011000000000";
        when 245 => y_in <= "10000000"; x_in <= "01110101"; z_correct<="1100010110000000";
        when 246 => y_in <= "10000000"; x_in <= "01110110"; z_correct<="1100010100000000";
        when 247 => y_in <= "10000000"; x_in <= "01110111"; z_correct<="1100010010000000";
        when 248 => y_in <= "10000000"; x_in <= "01111000"; z_correct<="1100010000000000";
        when 249 => y_in <= "10000000"; x_in <= "01111001"; z_correct<="1100001110000000";
        when 250 => y_in <= "10000000"; x_in <= "01111010"; z_correct<="1100001100000000";
        when 251 => y_in <= "10000000"; x_in <= "01111011"; z_correct<="1100001010000000";
        when 252 => y_in <= "10000000"; x_in <= "01111100"; z_correct<="1100001000000000";
        when 253 => y_in <= "10000000"; x_in <= "01111101"; z_correct<="1100000110000000";
        when 254 => y_in <= "10000000"; x_in <= "01111110"; z_correct<="1100000100000000";
        when 255 => y_in <= "10000000"; x_in <= "01111111"; z_correct<="1100000010000000";
        when 256 => y_in <= "10000001"; x_in <= "10000000"; z_correct<="0011111110000000";
        when 257 => y_in <= "10000001"; x_in <= "10000001"; z_correct<="0011111100000001";
        when 258 => y_in <= "10000001"; x_in <= "10000010"; z_correct<="0011111010000010";
        when 259 => y_in <= "10000001"; x_in <= "10000011"; z_correct<="0011111000000011";
        when 260 => y_in <= "10000001"; x_in <= "10000100"; z_correct<="0011110110000100";
        when 261 => y_in <= "10000001"; x_in <= "10000101"; z_correct<="0011110100000101";
        when 262 => y_in <= "10000001"; x_in <= "10000110"; z_correct<="0011110010000110";
        when 263 => y_in <= "10000001"; x_in <= "10000111"; z_correct<="0011110000000111";
        when 264 => y_in <= "10000001"; x_in <= "10001000"; z_correct<="0011101110001000";
        when 265 => y_in <= "10000001"; x_in <= "10001001"; z_correct<="0011101100001001";
        when 266 => y_in <= "10000001"; x_in <= "10001010"; z_correct<="0011101010001010";
        when 267 => y_in <= "10000001"; x_in <= "10001011"; z_correct<="0011101000001011";
        when 268 => y_in <= "10000001"; x_in <= "10001100"; z_correct<="0011100110001100";
        when 269 => y_in <= "10000001"; x_in <= "10001101"; z_correct<="0011100100001101";
        when 270 => y_in <= "10000001"; x_in <= "10001110"; z_correct<="0011100010001110";
        when 271 => y_in <= "10000001"; x_in <= "10001111"; z_correct<="0011100000001111";
        when 272 => y_in <= "10000001"; x_in <= "10010000"; z_correct<="0011011110010000";
        when 273 => y_in <= "10000001"; x_in <= "10010001"; z_correct<="0011011100010001";
        when 274 => y_in <= "10000001"; x_in <= "10010010"; z_correct<="0011011010010010";
        when 275 => y_in <= "10000001"; x_in <= "10010011"; z_correct<="0011011000010011";
        when 276 => y_in <= "10000001"; x_in <= "10010100"; z_correct<="0011010110010100";
        when 277 => y_in <= "10000001"; x_in <= "10010101"; z_correct<="0011010100010101";
        when 278 => y_in <= "10000001"; x_in <= "10010110"; z_correct<="0011010010010110";
        when 279 => y_in <= "10000001"; x_in <= "10010111"; z_correct<="0011010000010111";
        when 280 => y_in <= "10000001"; x_in <= "10011000"; z_correct<="0011001110011000";
        when 281 => y_in <= "10000001"; x_in <= "10011001"; z_correct<="0011001100011001";
        when 282 => y_in <= "10000001"; x_in <= "10011010"; z_correct<="0011001010011010";
        when 283 => y_in <= "10000001"; x_in <= "10011011"; z_correct<="0011001000011011";
        when 284 => y_in <= "10000001"; x_in <= "10011100"; z_correct<="0011000110011100";
        when 285 => y_in <= "10000001"; x_in <= "10011101"; z_correct<="0011000100011101";
        when 286 => y_in <= "10000001"; x_in <= "10011110"; z_correct<="0011000010011110";
        when 287 => y_in <= "10000001"; x_in <= "10011111"; z_correct<="0011000000011111";
        when 288 => y_in <= "10000001"; x_in <= "10100000"; z_correct<="0010111110100000";
        when 289 => y_in <= "10000001"; x_in <= "10100001"; z_correct<="0010111100100001";
        when 290 => y_in <= "10000001"; x_in <= "10100010"; z_correct<="0010111010100010";
        when 291 => y_in <= "10000001"; x_in <= "10100011"; z_correct<="0010111000100011";
        when 292 => y_in <= "10000001"; x_in <= "10100100"; z_correct<="0010110110100100";
        when 293 => y_in <= "10000001"; x_in <= "10100101"; z_correct<="0010110100100101";
        when 294 => y_in <= "10000001"; x_in <= "10100110"; z_correct<="0010110010100110";
        when 295 => y_in <= "10000001"; x_in <= "10100111"; z_correct<="0010110000100111";
        when 296 => y_in <= "10000001"; x_in <= "10101000"; z_correct<="0010101110101000";
        when 297 => y_in <= "10000001"; x_in <= "10101001"; z_correct<="0010101100101001";
        when 298 => y_in <= "10000001"; x_in <= "10101010"; z_correct<="0010101010101010";
        when 299 => y_in <= "10000001"; x_in <= "10101011"; z_correct<="0010101000101011";
        when 300 => y_in <= "10000001"; x_in <= "10101100"; z_correct<="0010100110101100";
        when 301 => y_in <= "10000001"; x_in <= "10101101"; z_correct<="0010100100101101";
        when 302 => y_in <= "10000001"; x_in <= "10101110"; z_correct<="0010100010101110";
        when 303 => y_in <= "10000001"; x_in <= "10101111"; z_correct<="0010100000101111";
        when 304 => y_in <= "10000001"; x_in <= "10110000"; z_correct<="0010011110110000";
        when 305 => y_in <= "10000001"; x_in <= "10110001"; z_correct<="0010011100110001";
        when 306 => y_in <= "10000001"; x_in <= "10110010"; z_correct<="0010011010110010";
        when 307 => y_in <= "10000001"; x_in <= "10110011"; z_correct<="0010011000110011";
        when 308 => y_in <= "10000001"; x_in <= "10110100"; z_correct<="0010010110110100";
        when 309 => y_in <= "10000001"; x_in <= "10110101"; z_correct<="0010010100110101";
        when 310 => y_in <= "10000001"; x_in <= "10110110"; z_correct<="0010010010110110";
        when 311 => y_in <= "10000001"; x_in <= "10110111"; z_correct<="0010010000110111";
        when 312 => y_in <= "10000001"; x_in <= "10111000"; z_correct<="0010001110111000";
        when 313 => y_in <= "10000001"; x_in <= "10111001"; z_correct<="0010001100111001";
        when 314 => y_in <= "10000001"; x_in <= "10111010"; z_correct<="0010001010111010";
        when 315 => y_in <= "10000001"; x_in <= "10111011"; z_correct<="0010001000111011";
        when 316 => y_in <= "10000001"; x_in <= "10111100"; z_correct<="0010000110111100";
        when 317 => y_in <= "10000001"; x_in <= "10111101"; z_correct<="0010000100111101";
        when 318 => y_in <= "10000001"; x_in <= "10111110"; z_correct<="0010000010111110";
        when 319 => y_in <= "10000001"; x_in <= "10111111"; z_correct<="0010000000111111";
        when 320 => y_in <= "10000001"; x_in <= "11000000"; z_correct<="0001111111000000";
        when 321 => y_in <= "10000001"; x_in <= "11000001"; z_correct<="0001111101000001";
        when 322 => y_in <= "10000001"; x_in <= "11000010"; z_correct<="0001111011000010";
        when 323 => y_in <= "10000001"; x_in <= "11000011"; z_correct<="0001111001000011";
        when 324 => y_in <= "10000001"; x_in <= "11000100"; z_correct<="0001110111000100";
        when 325 => y_in <= "10000001"; x_in <= "11000101"; z_correct<="0001110101000101";
        when 326 => y_in <= "10000001"; x_in <= "11000110"; z_correct<="0001110011000110";
        when 327 => y_in <= "10000001"; x_in <= "11000111"; z_correct<="0001110001000111";
        when 328 => y_in <= "10000001"; x_in <= "11001000"; z_correct<="0001101111001000";
        when 329 => y_in <= "10000001"; x_in <= "11001001"; z_correct<="0001101101001001";
        when 330 => y_in <= "10000001"; x_in <= "11001010"; z_correct<="0001101011001010";
        when 331 => y_in <= "10000001"; x_in <= "11001011"; z_correct<="0001101001001011";
        when 332 => y_in <= "10000001"; x_in <= "11001100"; z_correct<="0001100111001100";
        when 333 => y_in <= "10000001"; x_in <= "11001101"; z_correct<="0001100101001101";
        when 334 => y_in <= "10000001"; x_in <= "11001110"; z_correct<="0001100011001110";
        when 335 => y_in <= "10000001"; x_in <= "11001111"; z_correct<="0001100001001111";
        when 336 => y_in <= "10000001"; x_in <= "11010000"; z_correct<="0001011111010000";
        when 337 => y_in <= "10000001"; x_in <= "11010001"; z_correct<="0001011101010001";
        when 338 => y_in <= "10000001"; x_in <= "11010010"; z_correct<="0001011011010010";
        when 339 => y_in <= "10000001"; x_in <= "11010011"; z_correct<="0001011001010011";
        when 340 => y_in <= "10000001"; x_in <= "11010100"; z_correct<="0001010111010100";
        when 341 => y_in <= "10000001"; x_in <= "11010101"; z_correct<="0001010101010101";
        when 342 => y_in <= "10000001"; x_in <= "11010110"; z_correct<="0001010011010110";
        when 343 => y_in <= "10000001"; x_in <= "11010111"; z_correct<="0001010001010111";
        when 344 => y_in <= "10000001"; x_in <= "11011000"; z_correct<="0001001111011000";
        when 345 => y_in <= "10000001"; x_in <= "11011001"; z_correct<="0001001101011001";
        when 346 => y_in <= "10000001"; x_in <= "11011010"; z_correct<="0001001011011010";
        when 347 => y_in <= "10000001"; x_in <= "11011011"; z_correct<="0001001001011011";
        when 348 => y_in <= "10000001"; x_in <= "11011100"; z_correct<="0001000111011100";
        when 349 => y_in <= "10000001"; x_in <= "11011101"; z_correct<="0001000101011101";
        when 350 => y_in <= "10000001"; x_in <= "11011110"; z_correct<="0001000011011110";
        when 351 => y_in <= "10000001"; x_in <= "11011111"; z_correct<="0001000001011111";
        when 352 => y_in <= "10000001"; x_in <= "11100000"; z_correct<="0000111111100000";
        when 353 => y_in <= "10000001"; x_in <= "11100001"; z_correct<="0000111101100001";
        when 354 => y_in <= "10000001"; x_in <= "11100010"; z_correct<="0000111011100010";
        when 355 => y_in <= "10000001"; x_in <= "11100011"; z_correct<="0000111001100011";
        when 356 => y_in <= "10000001"; x_in <= "11100100"; z_correct<="0000110111100100";
        when 357 => y_in <= "10000001"; x_in <= "11100101"; z_correct<="0000110101100101";
        when 358 => y_in <= "10000001"; x_in <= "11100110"; z_correct<="0000110011100110";
        when 359 => y_in <= "10000001"; x_in <= "11100111"; z_correct<="0000110001100111";
        when 360 => y_in <= "10000001"; x_in <= "11101000"; z_correct<="0000101111101000";
        when 361 => y_in <= "10000001"; x_in <= "11101001"; z_correct<="0000101101101001";
        when 362 => y_in <= "10000001"; x_in <= "11101010"; z_correct<="0000101011101010";
        when 363 => y_in <= "10000001"; x_in <= "11101011"; z_correct<="0000101001101011";
        when 364 => y_in <= "10000001"; x_in <= "11101100"; z_correct<="0000100111101100";
        when 365 => y_in <= "10000001"; x_in <= "11101101"; z_correct<="0000100101101101";
        when 366 => y_in <= "10000001"; x_in <= "11101110"; z_correct<="0000100011101110";
        when 367 => y_in <= "10000001"; x_in <= "11101111"; z_correct<="0000100001101111";
        when 368 => y_in <= "10000001"; x_in <= "11110000"; z_correct<="0000011111110000";
        when 369 => y_in <= "10000001"; x_in <= "11110001"; z_correct<="0000011101110001";
        when 370 => y_in <= "10000001"; x_in <= "11110010"; z_correct<="0000011011110010";
        when 371 => y_in <= "10000001"; x_in <= "11110011"; z_correct<="0000011001110011";
        when 372 => y_in <= "10000001"; x_in <= "11110100"; z_correct<="0000010111110100";
        when 373 => y_in <= "10000001"; x_in <= "11110101"; z_correct<="0000010101110101";
        when 374 => y_in <= "10000001"; x_in <= "11110110"; z_correct<="0000010011110110";
        when 375 => y_in <= "10000001"; x_in <= "11110111"; z_correct<="0000010001110111";
        when 376 => y_in <= "10000001"; x_in <= "11111000"; z_correct<="0000001111111000";
        when 377 => y_in <= "10000001"; x_in <= "11111001"; z_correct<="0000001101111001";
        when 378 => y_in <= "10000001"; x_in <= "11111010"; z_correct<="0000001011111010";
        when 379 => y_in <= "10000001"; x_in <= "11111011"; z_correct<="0000001001111011";
        when 380 => y_in <= "10000001"; x_in <= "11111100"; z_correct<="0000000111111100";
        when 381 => y_in <= "10000001"; x_in <= "11111101"; z_correct<="0000000101111101";
        when 382 => y_in <= "10000001"; x_in <= "11111110"; z_correct<="0000000011111110";
        when 383 => y_in <= "10000001"; x_in <= "11111111"; z_correct<="0000000001111111";
        when 384 => y_in <= "10000001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 385 => y_in <= "10000001"; x_in <= "00000001"; z_correct<="1111111110000001";
        when 386 => y_in <= "10000001"; x_in <= "00000010"; z_correct<="1111111100000010";
        when 387 => y_in <= "10000001"; x_in <= "00000011"; z_correct<="1111111010000011";
        when 388 => y_in <= "10000001"; x_in <= "00000100"; z_correct<="1111111000000100";
        when 389 => y_in <= "10000001"; x_in <= "00000101"; z_correct<="1111110110000101";
        when 390 => y_in <= "10000001"; x_in <= "00000110"; z_correct<="1111110100000110";
        when 391 => y_in <= "10000001"; x_in <= "00000111"; z_correct<="1111110010000111";
        when 392 => y_in <= "10000001"; x_in <= "00001000"; z_correct<="1111110000001000";
        when 393 => y_in <= "10000001"; x_in <= "00001001"; z_correct<="1111101110001001";
        when 394 => y_in <= "10000001"; x_in <= "00001010"; z_correct<="1111101100001010";
        when 395 => y_in <= "10000001"; x_in <= "00001011"; z_correct<="1111101010001011";
        when 396 => y_in <= "10000001"; x_in <= "00001100"; z_correct<="1111101000001100";
        when 397 => y_in <= "10000001"; x_in <= "00001101"; z_correct<="1111100110001101";
        when 398 => y_in <= "10000001"; x_in <= "00001110"; z_correct<="1111100100001110";
        when 399 => y_in <= "10000001"; x_in <= "00001111"; z_correct<="1111100010001111";
        when 400 => y_in <= "10000001"; x_in <= "00010000"; z_correct<="1111100000010000";
        when 401 => y_in <= "10000001"; x_in <= "00010001"; z_correct<="1111011110010001";
        when 402 => y_in <= "10000001"; x_in <= "00010010"; z_correct<="1111011100010010";
        when 403 => y_in <= "10000001"; x_in <= "00010011"; z_correct<="1111011010010011";
        when 404 => y_in <= "10000001"; x_in <= "00010100"; z_correct<="1111011000010100";
        when 405 => y_in <= "10000001"; x_in <= "00010101"; z_correct<="1111010110010101";
        when 406 => y_in <= "10000001"; x_in <= "00010110"; z_correct<="1111010100010110";
        when 407 => y_in <= "10000001"; x_in <= "00010111"; z_correct<="1111010010010111";
        when 408 => y_in <= "10000001"; x_in <= "00011000"; z_correct<="1111010000011000";
        when 409 => y_in <= "10000001"; x_in <= "00011001"; z_correct<="1111001110011001";
        when 410 => y_in <= "10000001"; x_in <= "00011010"; z_correct<="1111001100011010";
        when 411 => y_in <= "10000001"; x_in <= "00011011"; z_correct<="1111001010011011";
        when 412 => y_in <= "10000001"; x_in <= "00011100"; z_correct<="1111001000011100";
        when 413 => y_in <= "10000001"; x_in <= "00011101"; z_correct<="1111000110011101";
        when 414 => y_in <= "10000001"; x_in <= "00011110"; z_correct<="1111000100011110";
        when 415 => y_in <= "10000001"; x_in <= "00011111"; z_correct<="1111000010011111";
        when 416 => y_in <= "10000001"; x_in <= "00100000"; z_correct<="1111000000100000";
        when 417 => y_in <= "10000001"; x_in <= "00100001"; z_correct<="1110111110100001";
        when 418 => y_in <= "10000001"; x_in <= "00100010"; z_correct<="1110111100100010";
        when 419 => y_in <= "10000001"; x_in <= "00100011"; z_correct<="1110111010100011";
        when 420 => y_in <= "10000001"; x_in <= "00100100"; z_correct<="1110111000100100";
        when 421 => y_in <= "10000001"; x_in <= "00100101"; z_correct<="1110110110100101";
        when 422 => y_in <= "10000001"; x_in <= "00100110"; z_correct<="1110110100100110";
        when 423 => y_in <= "10000001"; x_in <= "00100111"; z_correct<="1110110010100111";
        when 424 => y_in <= "10000001"; x_in <= "00101000"; z_correct<="1110110000101000";
        when 425 => y_in <= "10000001"; x_in <= "00101001"; z_correct<="1110101110101001";
        when 426 => y_in <= "10000001"; x_in <= "00101010"; z_correct<="1110101100101010";
        when 427 => y_in <= "10000001"; x_in <= "00101011"; z_correct<="1110101010101011";
        when 428 => y_in <= "10000001"; x_in <= "00101100"; z_correct<="1110101000101100";
        when 429 => y_in <= "10000001"; x_in <= "00101101"; z_correct<="1110100110101101";
        when 430 => y_in <= "10000001"; x_in <= "00101110"; z_correct<="1110100100101110";
        when 431 => y_in <= "10000001"; x_in <= "00101111"; z_correct<="1110100010101111";
        when 432 => y_in <= "10000001"; x_in <= "00110000"; z_correct<="1110100000110000";
        when 433 => y_in <= "10000001"; x_in <= "00110001"; z_correct<="1110011110110001";
        when 434 => y_in <= "10000001"; x_in <= "00110010"; z_correct<="1110011100110010";
        when 435 => y_in <= "10000001"; x_in <= "00110011"; z_correct<="1110011010110011";
        when 436 => y_in <= "10000001"; x_in <= "00110100"; z_correct<="1110011000110100";
        when 437 => y_in <= "10000001"; x_in <= "00110101"; z_correct<="1110010110110101";
        when 438 => y_in <= "10000001"; x_in <= "00110110"; z_correct<="1110010100110110";
        when 439 => y_in <= "10000001"; x_in <= "00110111"; z_correct<="1110010010110111";
        when 440 => y_in <= "10000001"; x_in <= "00111000"; z_correct<="1110010000111000";
        when 441 => y_in <= "10000001"; x_in <= "00111001"; z_correct<="1110001110111001";
        when 442 => y_in <= "10000001"; x_in <= "00111010"; z_correct<="1110001100111010";
        when 443 => y_in <= "10000001"; x_in <= "00111011"; z_correct<="1110001010111011";
        when 444 => y_in <= "10000001"; x_in <= "00111100"; z_correct<="1110001000111100";
        when 445 => y_in <= "10000001"; x_in <= "00111101"; z_correct<="1110000110111101";
        when 446 => y_in <= "10000001"; x_in <= "00111110"; z_correct<="1110000100111110";
        when 447 => y_in <= "10000001"; x_in <= "00111111"; z_correct<="1110000010111111";
        when 448 => y_in <= "10000001"; x_in <= "01000000"; z_correct<="1110000001000000";
        when 449 => y_in <= "10000001"; x_in <= "01000001"; z_correct<="1101111111000001";
        when 450 => y_in <= "10000001"; x_in <= "01000010"; z_correct<="1101111101000010";
        when 451 => y_in <= "10000001"; x_in <= "01000011"; z_correct<="1101111011000011";
        when 452 => y_in <= "10000001"; x_in <= "01000100"; z_correct<="1101111001000100";
        when 453 => y_in <= "10000001"; x_in <= "01000101"; z_correct<="1101110111000101";
        when 454 => y_in <= "10000001"; x_in <= "01000110"; z_correct<="1101110101000110";
        when 455 => y_in <= "10000001"; x_in <= "01000111"; z_correct<="1101110011000111";
        when 456 => y_in <= "10000001"; x_in <= "01001000"; z_correct<="1101110001001000";
        when 457 => y_in <= "10000001"; x_in <= "01001001"; z_correct<="1101101111001001";
        when 458 => y_in <= "10000001"; x_in <= "01001010"; z_correct<="1101101101001010";
        when 459 => y_in <= "10000001"; x_in <= "01001011"; z_correct<="1101101011001011";
        when 460 => y_in <= "10000001"; x_in <= "01001100"; z_correct<="1101101001001100";
        when 461 => y_in <= "10000001"; x_in <= "01001101"; z_correct<="1101100111001101";
        when 462 => y_in <= "10000001"; x_in <= "01001110"; z_correct<="1101100101001110";
        when 463 => y_in <= "10000001"; x_in <= "01001111"; z_correct<="1101100011001111";
        when 464 => y_in <= "10000001"; x_in <= "01010000"; z_correct<="1101100001010000";
        when 465 => y_in <= "10000001"; x_in <= "01010001"; z_correct<="1101011111010001";
        when 466 => y_in <= "10000001"; x_in <= "01010010"; z_correct<="1101011101010010";
        when 467 => y_in <= "10000001"; x_in <= "01010011"; z_correct<="1101011011010011";
        when 468 => y_in <= "10000001"; x_in <= "01010100"; z_correct<="1101011001010100";
        when 469 => y_in <= "10000001"; x_in <= "01010101"; z_correct<="1101010111010101";
        when 470 => y_in <= "10000001"; x_in <= "01010110"; z_correct<="1101010101010110";
        when 471 => y_in <= "10000001"; x_in <= "01010111"; z_correct<="1101010011010111";
        when 472 => y_in <= "10000001"; x_in <= "01011000"; z_correct<="1101010001011000";
        when 473 => y_in <= "10000001"; x_in <= "01011001"; z_correct<="1101001111011001";
        when 474 => y_in <= "10000001"; x_in <= "01011010"; z_correct<="1101001101011010";
        when 475 => y_in <= "10000001"; x_in <= "01011011"; z_correct<="1101001011011011";
        when 476 => y_in <= "10000001"; x_in <= "01011100"; z_correct<="1101001001011100";
        when 477 => y_in <= "10000001"; x_in <= "01011101"; z_correct<="1101000111011101";
        when 478 => y_in <= "10000001"; x_in <= "01011110"; z_correct<="1101000101011110";
        when 479 => y_in <= "10000001"; x_in <= "01011111"; z_correct<="1101000011011111";
        when 480 => y_in <= "10000001"; x_in <= "01100000"; z_correct<="1101000001100000";
        when 481 => y_in <= "10000001"; x_in <= "01100001"; z_correct<="1100111111100001";
        when 482 => y_in <= "10000001"; x_in <= "01100010"; z_correct<="1100111101100010";
        when 483 => y_in <= "10000001"; x_in <= "01100011"; z_correct<="1100111011100011";
        when 484 => y_in <= "10000001"; x_in <= "01100100"; z_correct<="1100111001100100";
        when 485 => y_in <= "10000001"; x_in <= "01100101"; z_correct<="1100110111100101";
        when 486 => y_in <= "10000001"; x_in <= "01100110"; z_correct<="1100110101100110";
        when 487 => y_in <= "10000001"; x_in <= "01100111"; z_correct<="1100110011100111";
        when 488 => y_in <= "10000001"; x_in <= "01101000"; z_correct<="1100110001101000";
        when 489 => y_in <= "10000001"; x_in <= "01101001"; z_correct<="1100101111101001";
        when 490 => y_in <= "10000001"; x_in <= "01101010"; z_correct<="1100101101101010";
        when 491 => y_in <= "10000001"; x_in <= "01101011"; z_correct<="1100101011101011";
        when 492 => y_in <= "10000001"; x_in <= "01101100"; z_correct<="1100101001101100";
        when 493 => y_in <= "10000001"; x_in <= "01101101"; z_correct<="1100100111101101";
        when 494 => y_in <= "10000001"; x_in <= "01101110"; z_correct<="1100100101101110";
        when 495 => y_in <= "10000001"; x_in <= "01101111"; z_correct<="1100100011101111";
        when 496 => y_in <= "10000001"; x_in <= "01110000"; z_correct<="1100100001110000";
        when 497 => y_in <= "10000001"; x_in <= "01110001"; z_correct<="1100011111110001";
        when 498 => y_in <= "10000001"; x_in <= "01110010"; z_correct<="1100011101110010";
        when 499 => y_in <= "10000001"; x_in <= "01110011"; z_correct<="1100011011110011";
        when 500 => y_in <= "10000001"; x_in <= "01110100"; z_correct<="1100011001110100";
        when 501 => y_in <= "10000001"; x_in <= "01110101"; z_correct<="1100010111110101";
        when 502 => y_in <= "10000001"; x_in <= "01110110"; z_correct<="1100010101110110";
        when 503 => y_in <= "10000001"; x_in <= "01110111"; z_correct<="1100010011110111";
        when 504 => y_in <= "10000001"; x_in <= "01111000"; z_correct<="1100010001111000";
        when 505 => y_in <= "10000001"; x_in <= "01111001"; z_correct<="1100001111111001";
        when 506 => y_in <= "10000001"; x_in <= "01111010"; z_correct<="1100001101111010";
        when 507 => y_in <= "10000001"; x_in <= "01111011"; z_correct<="1100001011111011";
        when 508 => y_in <= "10000001"; x_in <= "01111100"; z_correct<="1100001001111100";
        when 509 => y_in <= "10000001"; x_in <= "01111101"; z_correct<="1100000111111101";
        when 510 => y_in <= "10000001"; x_in <= "01111110"; z_correct<="1100000101111110";
        when 511 => y_in <= "10000001"; x_in <= "01111111"; z_correct<="1100000011111111";
        when 512 => y_in <= "10000010"; x_in <= "10000000"; z_correct<="0011111100000000";
        when 513 => y_in <= "10000010"; x_in <= "10000001"; z_correct<="0011111010000010";
        when 514 => y_in <= "10000010"; x_in <= "10000010"; z_correct<="0011111000000100";
        when 515 => y_in <= "10000010"; x_in <= "10000011"; z_correct<="0011110110000110";
        when 516 => y_in <= "10000010"; x_in <= "10000100"; z_correct<="0011110100001000";
        when 517 => y_in <= "10000010"; x_in <= "10000101"; z_correct<="0011110010001010";
        when 518 => y_in <= "10000010"; x_in <= "10000110"; z_correct<="0011110000001100";
        when 519 => y_in <= "10000010"; x_in <= "10000111"; z_correct<="0011101110001110";
        when 520 => y_in <= "10000010"; x_in <= "10001000"; z_correct<="0011101100010000";
        when 521 => y_in <= "10000010"; x_in <= "10001001"; z_correct<="0011101010010010";
        when 522 => y_in <= "10000010"; x_in <= "10001010"; z_correct<="0011101000010100";
        when 523 => y_in <= "10000010"; x_in <= "10001011"; z_correct<="0011100110010110";
        when 524 => y_in <= "10000010"; x_in <= "10001100"; z_correct<="0011100100011000";
        when 525 => y_in <= "10000010"; x_in <= "10001101"; z_correct<="0011100010011010";
        when 526 => y_in <= "10000010"; x_in <= "10001110"; z_correct<="0011100000011100";
        when 527 => y_in <= "10000010"; x_in <= "10001111"; z_correct<="0011011110011110";
        when 528 => y_in <= "10000010"; x_in <= "10010000"; z_correct<="0011011100100000";
        when 529 => y_in <= "10000010"; x_in <= "10010001"; z_correct<="0011011010100010";
        when 530 => y_in <= "10000010"; x_in <= "10010010"; z_correct<="0011011000100100";
        when 531 => y_in <= "10000010"; x_in <= "10010011"; z_correct<="0011010110100110";
        when 532 => y_in <= "10000010"; x_in <= "10010100"; z_correct<="0011010100101000";
        when 533 => y_in <= "10000010"; x_in <= "10010101"; z_correct<="0011010010101010";
        when 534 => y_in <= "10000010"; x_in <= "10010110"; z_correct<="0011010000101100";
        when 535 => y_in <= "10000010"; x_in <= "10010111"; z_correct<="0011001110101110";
        when 536 => y_in <= "10000010"; x_in <= "10011000"; z_correct<="0011001100110000";
        when 537 => y_in <= "10000010"; x_in <= "10011001"; z_correct<="0011001010110010";
        when 538 => y_in <= "10000010"; x_in <= "10011010"; z_correct<="0011001000110100";
        when 539 => y_in <= "10000010"; x_in <= "10011011"; z_correct<="0011000110110110";
        when 540 => y_in <= "10000010"; x_in <= "10011100"; z_correct<="0011000100111000";
        when 541 => y_in <= "10000010"; x_in <= "10011101"; z_correct<="0011000010111010";
        when 542 => y_in <= "10000010"; x_in <= "10011110"; z_correct<="0011000000111100";
        when 543 => y_in <= "10000010"; x_in <= "10011111"; z_correct<="0010111110111110";
        when 544 => y_in <= "10000010"; x_in <= "10100000"; z_correct<="0010111101000000";
        when 545 => y_in <= "10000010"; x_in <= "10100001"; z_correct<="0010111011000010";
        when 546 => y_in <= "10000010"; x_in <= "10100010"; z_correct<="0010111001000100";
        when 547 => y_in <= "10000010"; x_in <= "10100011"; z_correct<="0010110111000110";
        when 548 => y_in <= "10000010"; x_in <= "10100100"; z_correct<="0010110101001000";
        when 549 => y_in <= "10000010"; x_in <= "10100101"; z_correct<="0010110011001010";
        when 550 => y_in <= "10000010"; x_in <= "10100110"; z_correct<="0010110001001100";
        when 551 => y_in <= "10000010"; x_in <= "10100111"; z_correct<="0010101111001110";
        when 552 => y_in <= "10000010"; x_in <= "10101000"; z_correct<="0010101101010000";
        when 553 => y_in <= "10000010"; x_in <= "10101001"; z_correct<="0010101011010010";
        when 554 => y_in <= "10000010"; x_in <= "10101010"; z_correct<="0010101001010100";
        when 555 => y_in <= "10000010"; x_in <= "10101011"; z_correct<="0010100111010110";
        when 556 => y_in <= "10000010"; x_in <= "10101100"; z_correct<="0010100101011000";
        when 557 => y_in <= "10000010"; x_in <= "10101101"; z_correct<="0010100011011010";
        when 558 => y_in <= "10000010"; x_in <= "10101110"; z_correct<="0010100001011100";
        when 559 => y_in <= "10000010"; x_in <= "10101111"; z_correct<="0010011111011110";
        when 560 => y_in <= "10000010"; x_in <= "10110000"; z_correct<="0010011101100000";
        when 561 => y_in <= "10000010"; x_in <= "10110001"; z_correct<="0010011011100010";
        when 562 => y_in <= "10000010"; x_in <= "10110010"; z_correct<="0010011001100100";
        when 563 => y_in <= "10000010"; x_in <= "10110011"; z_correct<="0010010111100110";
        when 564 => y_in <= "10000010"; x_in <= "10110100"; z_correct<="0010010101101000";
        when 565 => y_in <= "10000010"; x_in <= "10110101"; z_correct<="0010010011101010";
        when 566 => y_in <= "10000010"; x_in <= "10110110"; z_correct<="0010010001101100";
        when 567 => y_in <= "10000010"; x_in <= "10110111"; z_correct<="0010001111101110";
        when 568 => y_in <= "10000010"; x_in <= "10111000"; z_correct<="0010001101110000";
        when 569 => y_in <= "10000010"; x_in <= "10111001"; z_correct<="0010001011110010";
        when 570 => y_in <= "10000010"; x_in <= "10111010"; z_correct<="0010001001110100";
        when 571 => y_in <= "10000010"; x_in <= "10111011"; z_correct<="0010000111110110";
        when 572 => y_in <= "10000010"; x_in <= "10111100"; z_correct<="0010000101111000";
        when 573 => y_in <= "10000010"; x_in <= "10111101"; z_correct<="0010000011111010";
        when 574 => y_in <= "10000010"; x_in <= "10111110"; z_correct<="0010000001111100";
        when 575 => y_in <= "10000010"; x_in <= "10111111"; z_correct<="0001111111111110";
        when 576 => y_in <= "10000010"; x_in <= "11000000"; z_correct<="0001111110000000";
        when 577 => y_in <= "10000010"; x_in <= "11000001"; z_correct<="0001111100000010";
        when 578 => y_in <= "10000010"; x_in <= "11000010"; z_correct<="0001111010000100";
        when 579 => y_in <= "10000010"; x_in <= "11000011"; z_correct<="0001111000000110";
        when 580 => y_in <= "10000010"; x_in <= "11000100"; z_correct<="0001110110001000";
        when 581 => y_in <= "10000010"; x_in <= "11000101"; z_correct<="0001110100001010";
        when 582 => y_in <= "10000010"; x_in <= "11000110"; z_correct<="0001110010001100";
        when 583 => y_in <= "10000010"; x_in <= "11000111"; z_correct<="0001110000001110";
        when 584 => y_in <= "10000010"; x_in <= "11001000"; z_correct<="0001101110010000";
        when 585 => y_in <= "10000010"; x_in <= "11001001"; z_correct<="0001101100010010";
        when 586 => y_in <= "10000010"; x_in <= "11001010"; z_correct<="0001101010010100";
        when 587 => y_in <= "10000010"; x_in <= "11001011"; z_correct<="0001101000010110";
        when 588 => y_in <= "10000010"; x_in <= "11001100"; z_correct<="0001100110011000";
        when 589 => y_in <= "10000010"; x_in <= "11001101"; z_correct<="0001100100011010";
        when 590 => y_in <= "10000010"; x_in <= "11001110"; z_correct<="0001100010011100";
        when 591 => y_in <= "10000010"; x_in <= "11001111"; z_correct<="0001100000011110";
        when 592 => y_in <= "10000010"; x_in <= "11010000"; z_correct<="0001011110100000";
        when 593 => y_in <= "10000010"; x_in <= "11010001"; z_correct<="0001011100100010";
        when 594 => y_in <= "10000010"; x_in <= "11010010"; z_correct<="0001011010100100";
        when 595 => y_in <= "10000010"; x_in <= "11010011"; z_correct<="0001011000100110";
        when 596 => y_in <= "10000010"; x_in <= "11010100"; z_correct<="0001010110101000";
        when 597 => y_in <= "10000010"; x_in <= "11010101"; z_correct<="0001010100101010";
        when 598 => y_in <= "10000010"; x_in <= "11010110"; z_correct<="0001010010101100";
        when 599 => y_in <= "10000010"; x_in <= "11010111"; z_correct<="0001010000101110";
        when 600 => y_in <= "10000010"; x_in <= "11011000"; z_correct<="0001001110110000";
        when 601 => y_in <= "10000010"; x_in <= "11011001"; z_correct<="0001001100110010";
        when 602 => y_in <= "10000010"; x_in <= "11011010"; z_correct<="0001001010110100";
        when 603 => y_in <= "10000010"; x_in <= "11011011"; z_correct<="0001001000110110";
        when 604 => y_in <= "10000010"; x_in <= "11011100"; z_correct<="0001000110111000";
        when 605 => y_in <= "10000010"; x_in <= "11011101"; z_correct<="0001000100111010";
        when 606 => y_in <= "10000010"; x_in <= "11011110"; z_correct<="0001000010111100";
        when 607 => y_in <= "10000010"; x_in <= "11011111"; z_correct<="0001000000111110";
        when 608 => y_in <= "10000010"; x_in <= "11100000"; z_correct<="0000111111000000";
        when 609 => y_in <= "10000010"; x_in <= "11100001"; z_correct<="0000111101000010";
        when 610 => y_in <= "10000010"; x_in <= "11100010"; z_correct<="0000111011000100";
        when 611 => y_in <= "10000010"; x_in <= "11100011"; z_correct<="0000111001000110";
        when 612 => y_in <= "10000010"; x_in <= "11100100"; z_correct<="0000110111001000";
        when 613 => y_in <= "10000010"; x_in <= "11100101"; z_correct<="0000110101001010";
        when 614 => y_in <= "10000010"; x_in <= "11100110"; z_correct<="0000110011001100";
        when 615 => y_in <= "10000010"; x_in <= "11100111"; z_correct<="0000110001001110";
        when 616 => y_in <= "10000010"; x_in <= "11101000"; z_correct<="0000101111010000";
        when 617 => y_in <= "10000010"; x_in <= "11101001"; z_correct<="0000101101010010";
        when 618 => y_in <= "10000010"; x_in <= "11101010"; z_correct<="0000101011010100";
        when 619 => y_in <= "10000010"; x_in <= "11101011"; z_correct<="0000101001010110";
        when 620 => y_in <= "10000010"; x_in <= "11101100"; z_correct<="0000100111011000";
        when 621 => y_in <= "10000010"; x_in <= "11101101"; z_correct<="0000100101011010";
        when 622 => y_in <= "10000010"; x_in <= "11101110"; z_correct<="0000100011011100";
        when 623 => y_in <= "10000010"; x_in <= "11101111"; z_correct<="0000100001011110";
        when 624 => y_in <= "10000010"; x_in <= "11110000"; z_correct<="0000011111100000";
        when 625 => y_in <= "10000010"; x_in <= "11110001"; z_correct<="0000011101100010";
        when 626 => y_in <= "10000010"; x_in <= "11110010"; z_correct<="0000011011100100";
        when 627 => y_in <= "10000010"; x_in <= "11110011"; z_correct<="0000011001100110";
        when 628 => y_in <= "10000010"; x_in <= "11110100"; z_correct<="0000010111101000";
        when 629 => y_in <= "10000010"; x_in <= "11110101"; z_correct<="0000010101101010";
        when 630 => y_in <= "10000010"; x_in <= "11110110"; z_correct<="0000010011101100";
        when 631 => y_in <= "10000010"; x_in <= "11110111"; z_correct<="0000010001101110";
        when 632 => y_in <= "10000010"; x_in <= "11111000"; z_correct<="0000001111110000";
        when 633 => y_in <= "10000010"; x_in <= "11111001"; z_correct<="0000001101110010";
        when 634 => y_in <= "10000010"; x_in <= "11111010"; z_correct<="0000001011110100";
        when 635 => y_in <= "10000010"; x_in <= "11111011"; z_correct<="0000001001110110";
        when 636 => y_in <= "10000010"; x_in <= "11111100"; z_correct<="0000000111111000";
        when 637 => y_in <= "10000010"; x_in <= "11111101"; z_correct<="0000000101111010";
        when 638 => y_in <= "10000010"; x_in <= "11111110"; z_correct<="0000000011111100";
        when 639 => y_in <= "10000010"; x_in <= "11111111"; z_correct<="0000000001111110";
        when 640 => y_in <= "10000010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 641 => y_in <= "10000010"; x_in <= "00000001"; z_correct<="1111111110000010";
        when 642 => y_in <= "10000010"; x_in <= "00000010"; z_correct<="1111111100000100";
        when 643 => y_in <= "10000010"; x_in <= "00000011"; z_correct<="1111111010000110";
        when 644 => y_in <= "10000010"; x_in <= "00000100"; z_correct<="1111111000001000";
        when 645 => y_in <= "10000010"; x_in <= "00000101"; z_correct<="1111110110001010";
        when 646 => y_in <= "10000010"; x_in <= "00000110"; z_correct<="1111110100001100";
        when 647 => y_in <= "10000010"; x_in <= "00000111"; z_correct<="1111110010001110";
        when 648 => y_in <= "10000010"; x_in <= "00001000"; z_correct<="1111110000010000";
        when 649 => y_in <= "10000010"; x_in <= "00001001"; z_correct<="1111101110010010";
        when 650 => y_in <= "10000010"; x_in <= "00001010"; z_correct<="1111101100010100";
        when 651 => y_in <= "10000010"; x_in <= "00001011"; z_correct<="1111101010010110";
        when 652 => y_in <= "10000010"; x_in <= "00001100"; z_correct<="1111101000011000";
        when 653 => y_in <= "10000010"; x_in <= "00001101"; z_correct<="1111100110011010";
        when 654 => y_in <= "10000010"; x_in <= "00001110"; z_correct<="1111100100011100";
        when 655 => y_in <= "10000010"; x_in <= "00001111"; z_correct<="1111100010011110";
        when 656 => y_in <= "10000010"; x_in <= "00010000"; z_correct<="1111100000100000";
        when 657 => y_in <= "10000010"; x_in <= "00010001"; z_correct<="1111011110100010";
        when 658 => y_in <= "10000010"; x_in <= "00010010"; z_correct<="1111011100100100";
        when 659 => y_in <= "10000010"; x_in <= "00010011"; z_correct<="1111011010100110";
        when 660 => y_in <= "10000010"; x_in <= "00010100"; z_correct<="1111011000101000";
        when 661 => y_in <= "10000010"; x_in <= "00010101"; z_correct<="1111010110101010";
        when 662 => y_in <= "10000010"; x_in <= "00010110"; z_correct<="1111010100101100";
        when 663 => y_in <= "10000010"; x_in <= "00010111"; z_correct<="1111010010101110";
        when 664 => y_in <= "10000010"; x_in <= "00011000"; z_correct<="1111010000110000";
        when 665 => y_in <= "10000010"; x_in <= "00011001"; z_correct<="1111001110110010";
        when 666 => y_in <= "10000010"; x_in <= "00011010"; z_correct<="1111001100110100";
        when 667 => y_in <= "10000010"; x_in <= "00011011"; z_correct<="1111001010110110";
        when 668 => y_in <= "10000010"; x_in <= "00011100"; z_correct<="1111001000111000";
        when 669 => y_in <= "10000010"; x_in <= "00011101"; z_correct<="1111000110111010";
        when 670 => y_in <= "10000010"; x_in <= "00011110"; z_correct<="1111000100111100";
        when 671 => y_in <= "10000010"; x_in <= "00011111"; z_correct<="1111000010111110";
        when 672 => y_in <= "10000010"; x_in <= "00100000"; z_correct<="1111000001000000";
        when 673 => y_in <= "10000010"; x_in <= "00100001"; z_correct<="1110111111000010";
        when 674 => y_in <= "10000010"; x_in <= "00100010"; z_correct<="1110111101000100";
        when 675 => y_in <= "10000010"; x_in <= "00100011"; z_correct<="1110111011000110";
        when 676 => y_in <= "10000010"; x_in <= "00100100"; z_correct<="1110111001001000";
        when 677 => y_in <= "10000010"; x_in <= "00100101"; z_correct<="1110110111001010";
        when 678 => y_in <= "10000010"; x_in <= "00100110"; z_correct<="1110110101001100";
        when 679 => y_in <= "10000010"; x_in <= "00100111"; z_correct<="1110110011001110";
        when 680 => y_in <= "10000010"; x_in <= "00101000"; z_correct<="1110110001010000";
        when 681 => y_in <= "10000010"; x_in <= "00101001"; z_correct<="1110101111010010";
        when 682 => y_in <= "10000010"; x_in <= "00101010"; z_correct<="1110101101010100";
        when 683 => y_in <= "10000010"; x_in <= "00101011"; z_correct<="1110101011010110";
        when 684 => y_in <= "10000010"; x_in <= "00101100"; z_correct<="1110101001011000";
        when 685 => y_in <= "10000010"; x_in <= "00101101"; z_correct<="1110100111011010";
        when 686 => y_in <= "10000010"; x_in <= "00101110"; z_correct<="1110100101011100";
        when 687 => y_in <= "10000010"; x_in <= "00101111"; z_correct<="1110100011011110";
        when 688 => y_in <= "10000010"; x_in <= "00110000"; z_correct<="1110100001100000";
        when 689 => y_in <= "10000010"; x_in <= "00110001"; z_correct<="1110011111100010";
        when 690 => y_in <= "10000010"; x_in <= "00110010"; z_correct<="1110011101100100";
        when 691 => y_in <= "10000010"; x_in <= "00110011"; z_correct<="1110011011100110";
        when 692 => y_in <= "10000010"; x_in <= "00110100"; z_correct<="1110011001101000";
        when 693 => y_in <= "10000010"; x_in <= "00110101"; z_correct<="1110010111101010";
        when 694 => y_in <= "10000010"; x_in <= "00110110"; z_correct<="1110010101101100";
        when 695 => y_in <= "10000010"; x_in <= "00110111"; z_correct<="1110010011101110";
        when 696 => y_in <= "10000010"; x_in <= "00111000"; z_correct<="1110010001110000";
        when 697 => y_in <= "10000010"; x_in <= "00111001"; z_correct<="1110001111110010";
        when 698 => y_in <= "10000010"; x_in <= "00111010"; z_correct<="1110001101110100";
        when 699 => y_in <= "10000010"; x_in <= "00111011"; z_correct<="1110001011110110";
        when 700 => y_in <= "10000010"; x_in <= "00111100"; z_correct<="1110001001111000";
        when 701 => y_in <= "10000010"; x_in <= "00111101"; z_correct<="1110000111111010";
        when 702 => y_in <= "10000010"; x_in <= "00111110"; z_correct<="1110000101111100";
        when 703 => y_in <= "10000010"; x_in <= "00111111"; z_correct<="1110000011111110";
        when 704 => y_in <= "10000010"; x_in <= "01000000"; z_correct<="1110000010000000";
        when 705 => y_in <= "10000010"; x_in <= "01000001"; z_correct<="1110000000000010";
        when 706 => y_in <= "10000010"; x_in <= "01000010"; z_correct<="1101111110000100";
        when 707 => y_in <= "10000010"; x_in <= "01000011"; z_correct<="1101111100000110";
        when 708 => y_in <= "10000010"; x_in <= "01000100"; z_correct<="1101111010001000";
        when 709 => y_in <= "10000010"; x_in <= "01000101"; z_correct<="1101111000001010";
        when 710 => y_in <= "10000010"; x_in <= "01000110"; z_correct<="1101110110001100";
        when 711 => y_in <= "10000010"; x_in <= "01000111"; z_correct<="1101110100001110";
        when 712 => y_in <= "10000010"; x_in <= "01001000"; z_correct<="1101110010010000";
        when 713 => y_in <= "10000010"; x_in <= "01001001"; z_correct<="1101110000010010";
        when 714 => y_in <= "10000010"; x_in <= "01001010"; z_correct<="1101101110010100";
        when 715 => y_in <= "10000010"; x_in <= "01001011"; z_correct<="1101101100010110";
        when 716 => y_in <= "10000010"; x_in <= "01001100"; z_correct<="1101101010011000";
        when 717 => y_in <= "10000010"; x_in <= "01001101"; z_correct<="1101101000011010";
        when 718 => y_in <= "10000010"; x_in <= "01001110"; z_correct<="1101100110011100";
        when 719 => y_in <= "10000010"; x_in <= "01001111"; z_correct<="1101100100011110";
        when 720 => y_in <= "10000010"; x_in <= "01010000"; z_correct<="1101100010100000";
        when 721 => y_in <= "10000010"; x_in <= "01010001"; z_correct<="1101100000100010";
        when 722 => y_in <= "10000010"; x_in <= "01010010"; z_correct<="1101011110100100";
        when 723 => y_in <= "10000010"; x_in <= "01010011"; z_correct<="1101011100100110";
        when 724 => y_in <= "10000010"; x_in <= "01010100"; z_correct<="1101011010101000";
        when 725 => y_in <= "10000010"; x_in <= "01010101"; z_correct<="1101011000101010";
        when 726 => y_in <= "10000010"; x_in <= "01010110"; z_correct<="1101010110101100";
        when 727 => y_in <= "10000010"; x_in <= "01010111"; z_correct<="1101010100101110";
        when 728 => y_in <= "10000010"; x_in <= "01011000"; z_correct<="1101010010110000";
        when 729 => y_in <= "10000010"; x_in <= "01011001"; z_correct<="1101010000110010";
        when 730 => y_in <= "10000010"; x_in <= "01011010"; z_correct<="1101001110110100";
        when 731 => y_in <= "10000010"; x_in <= "01011011"; z_correct<="1101001100110110";
        when 732 => y_in <= "10000010"; x_in <= "01011100"; z_correct<="1101001010111000";
        when 733 => y_in <= "10000010"; x_in <= "01011101"; z_correct<="1101001000111010";
        when 734 => y_in <= "10000010"; x_in <= "01011110"; z_correct<="1101000110111100";
        when 735 => y_in <= "10000010"; x_in <= "01011111"; z_correct<="1101000100111110";
        when 736 => y_in <= "10000010"; x_in <= "01100000"; z_correct<="1101000011000000";
        when 737 => y_in <= "10000010"; x_in <= "01100001"; z_correct<="1101000001000010";
        when 738 => y_in <= "10000010"; x_in <= "01100010"; z_correct<="1100111111000100";
        when 739 => y_in <= "10000010"; x_in <= "01100011"; z_correct<="1100111101000110";
        when 740 => y_in <= "10000010"; x_in <= "01100100"; z_correct<="1100111011001000";
        when 741 => y_in <= "10000010"; x_in <= "01100101"; z_correct<="1100111001001010";
        when 742 => y_in <= "10000010"; x_in <= "01100110"; z_correct<="1100110111001100";
        when 743 => y_in <= "10000010"; x_in <= "01100111"; z_correct<="1100110101001110";
        when 744 => y_in <= "10000010"; x_in <= "01101000"; z_correct<="1100110011010000";
        when 745 => y_in <= "10000010"; x_in <= "01101001"; z_correct<="1100110001010010";
        when 746 => y_in <= "10000010"; x_in <= "01101010"; z_correct<="1100101111010100";
        when 747 => y_in <= "10000010"; x_in <= "01101011"; z_correct<="1100101101010110";
        when 748 => y_in <= "10000010"; x_in <= "01101100"; z_correct<="1100101011011000";
        when 749 => y_in <= "10000010"; x_in <= "01101101"; z_correct<="1100101001011010";
        when 750 => y_in <= "10000010"; x_in <= "01101110"; z_correct<="1100100111011100";
        when 751 => y_in <= "10000010"; x_in <= "01101111"; z_correct<="1100100101011110";
        when 752 => y_in <= "10000010"; x_in <= "01110000"; z_correct<="1100100011100000";
        when 753 => y_in <= "10000010"; x_in <= "01110001"; z_correct<="1100100001100010";
        when 754 => y_in <= "10000010"; x_in <= "01110010"; z_correct<="1100011111100100";
        when 755 => y_in <= "10000010"; x_in <= "01110011"; z_correct<="1100011101100110";
        when 756 => y_in <= "10000010"; x_in <= "01110100"; z_correct<="1100011011101000";
        when 757 => y_in <= "10000010"; x_in <= "01110101"; z_correct<="1100011001101010";
        when 758 => y_in <= "10000010"; x_in <= "01110110"; z_correct<="1100010111101100";
        when 759 => y_in <= "10000010"; x_in <= "01110111"; z_correct<="1100010101101110";
        when 760 => y_in <= "10000010"; x_in <= "01111000"; z_correct<="1100010011110000";
        when 761 => y_in <= "10000010"; x_in <= "01111001"; z_correct<="1100010001110010";
        when 762 => y_in <= "10000010"; x_in <= "01111010"; z_correct<="1100001111110100";
        when 763 => y_in <= "10000010"; x_in <= "01111011"; z_correct<="1100001101110110";
        when 764 => y_in <= "10000010"; x_in <= "01111100"; z_correct<="1100001011111000";
        when 765 => y_in <= "10000010"; x_in <= "01111101"; z_correct<="1100001001111010";
        when 766 => y_in <= "10000010"; x_in <= "01111110"; z_correct<="1100000111111100";
        when 767 => y_in <= "10000010"; x_in <= "01111111"; z_correct<="1100000101111110";
        when 768 => y_in <= "10000011"; x_in <= "10000000"; z_correct<="0011111010000000";
        when 769 => y_in <= "10000011"; x_in <= "10000001"; z_correct<="0011111000000011";
        when 770 => y_in <= "10000011"; x_in <= "10000010"; z_correct<="0011110110000110";
        when 771 => y_in <= "10000011"; x_in <= "10000011"; z_correct<="0011110100001001";
        when 772 => y_in <= "10000011"; x_in <= "10000100"; z_correct<="0011110010001100";
        when 773 => y_in <= "10000011"; x_in <= "10000101"; z_correct<="0011110000001111";
        when 774 => y_in <= "10000011"; x_in <= "10000110"; z_correct<="0011101110010010";
        when 775 => y_in <= "10000011"; x_in <= "10000111"; z_correct<="0011101100010101";
        when 776 => y_in <= "10000011"; x_in <= "10001000"; z_correct<="0011101010011000";
        when 777 => y_in <= "10000011"; x_in <= "10001001"; z_correct<="0011101000011011";
        when 778 => y_in <= "10000011"; x_in <= "10001010"; z_correct<="0011100110011110";
        when 779 => y_in <= "10000011"; x_in <= "10001011"; z_correct<="0011100100100001";
        when 780 => y_in <= "10000011"; x_in <= "10001100"; z_correct<="0011100010100100";
        when 781 => y_in <= "10000011"; x_in <= "10001101"; z_correct<="0011100000100111";
        when 782 => y_in <= "10000011"; x_in <= "10001110"; z_correct<="0011011110101010";
        when 783 => y_in <= "10000011"; x_in <= "10001111"; z_correct<="0011011100101101";
        when 784 => y_in <= "10000011"; x_in <= "10010000"; z_correct<="0011011010110000";
        when 785 => y_in <= "10000011"; x_in <= "10010001"; z_correct<="0011011000110011";
        when 786 => y_in <= "10000011"; x_in <= "10010010"; z_correct<="0011010110110110";
        when 787 => y_in <= "10000011"; x_in <= "10010011"; z_correct<="0011010100111001";
        when 788 => y_in <= "10000011"; x_in <= "10010100"; z_correct<="0011010010111100";
        when 789 => y_in <= "10000011"; x_in <= "10010101"; z_correct<="0011010000111111";
        when 790 => y_in <= "10000011"; x_in <= "10010110"; z_correct<="0011001111000010";
        when 791 => y_in <= "10000011"; x_in <= "10010111"; z_correct<="0011001101000101";
        when 792 => y_in <= "10000011"; x_in <= "10011000"; z_correct<="0011001011001000";
        when 793 => y_in <= "10000011"; x_in <= "10011001"; z_correct<="0011001001001011";
        when 794 => y_in <= "10000011"; x_in <= "10011010"; z_correct<="0011000111001110";
        when 795 => y_in <= "10000011"; x_in <= "10011011"; z_correct<="0011000101010001";
        when 796 => y_in <= "10000011"; x_in <= "10011100"; z_correct<="0011000011010100";
        when 797 => y_in <= "10000011"; x_in <= "10011101"; z_correct<="0011000001010111";
        when 798 => y_in <= "10000011"; x_in <= "10011110"; z_correct<="0010111111011010";
        when 799 => y_in <= "10000011"; x_in <= "10011111"; z_correct<="0010111101011101";
        when 800 => y_in <= "10000011"; x_in <= "10100000"; z_correct<="0010111011100000";
        when 801 => y_in <= "10000011"; x_in <= "10100001"; z_correct<="0010111001100011";
        when 802 => y_in <= "10000011"; x_in <= "10100010"; z_correct<="0010110111100110";
        when 803 => y_in <= "10000011"; x_in <= "10100011"; z_correct<="0010110101101001";
        when 804 => y_in <= "10000011"; x_in <= "10100100"; z_correct<="0010110011101100";
        when 805 => y_in <= "10000011"; x_in <= "10100101"; z_correct<="0010110001101111";
        when 806 => y_in <= "10000011"; x_in <= "10100110"; z_correct<="0010101111110010";
        when 807 => y_in <= "10000011"; x_in <= "10100111"; z_correct<="0010101101110101";
        when 808 => y_in <= "10000011"; x_in <= "10101000"; z_correct<="0010101011111000";
        when 809 => y_in <= "10000011"; x_in <= "10101001"; z_correct<="0010101001111011";
        when 810 => y_in <= "10000011"; x_in <= "10101010"; z_correct<="0010100111111110";
        when 811 => y_in <= "10000011"; x_in <= "10101011"; z_correct<="0010100110000001";
        when 812 => y_in <= "10000011"; x_in <= "10101100"; z_correct<="0010100100000100";
        when 813 => y_in <= "10000011"; x_in <= "10101101"; z_correct<="0010100010000111";
        when 814 => y_in <= "10000011"; x_in <= "10101110"; z_correct<="0010100000001010";
        when 815 => y_in <= "10000011"; x_in <= "10101111"; z_correct<="0010011110001101";
        when 816 => y_in <= "10000011"; x_in <= "10110000"; z_correct<="0010011100010000";
        when 817 => y_in <= "10000011"; x_in <= "10110001"; z_correct<="0010011010010011";
        when 818 => y_in <= "10000011"; x_in <= "10110010"; z_correct<="0010011000010110";
        when 819 => y_in <= "10000011"; x_in <= "10110011"; z_correct<="0010010110011001";
        when 820 => y_in <= "10000011"; x_in <= "10110100"; z_correct<="0010010100011100";
        when 821 => y_in <= "10000011"; x_in <= "10110101"; z_correct<="0010010010011111";
        when 822 => y_in <= "10000011"; x_in <= "10110110"; z_correct<="0010010000100010";
        when 823 => y_in <= "10000011"; x_in <= "10110111"; z_correct<="0010001110100101";
        when 824 => y_in <= "10000011"; x_in <= "10111000"; z_correct<="0010001100101000";
        when 825 => y_in <= "10000011"; x_in <= "10111001"; z_correct<="0010001010101011";
        when 826 => y_in <= "10000011"; x_in <= "10111010"; z_correct<="0010001000101110";
        when 827 => y_in <= "10000011"; x_in <= "10111011"; z_correct<="0010000110110001";
        when 828 => y_in <= "10000011"; x_in <= "10111100"; z_correct<="0010000100110100";
        when 829 => y_in <= "10000011"; x_in <= "10111101"; z_correct<="0010000010110111";
        when 830 => y_in <= "10000011"; x_in <= "10111110"; z_correct<="0010000000111010";
        when 831 => y_in <= "10000011"; x_in <= "10111111"; z_correct<="0001111110111101";
        when 832 => y_in <= "10000011"; x_in <= "11000000"; z_correct<="0001111101000000";
        when 833 => y_in <= "10000011"; x_in <= "11000001"; z_correct<="0001111011000011";
        when 834 => y_in <= "10000011"; x_in <= "11000010"; z_correct<="0001111001000110";
        when 835 => y_in <= "10000011"; x_in <= "11000011"; z_correct<="0001110111001001";
        when 836 => y_in <= "10000011"; x_in <= "11000100"; z_correct<="0001110101001100";
        when 837 => y_in <= "10000011"; x_in <= "11000101"; z_correct<="0001110011001111";
        when 838 => y_in <= "10000011"; x_in <= "11000110"; z_correct<="0001110001010010";
        when 839 => y_in <= "10000011"; x_in <= "11000111"; z_correct<="0001101111010101";
        when 840 => y_in <= "10000011"; x_in <= "11001000"; z_correct<="0001101101011000";
        when 841 => y_in <= "10000011"; x_in <= "11001001"; z_correct<="0001101011011011";
        when 842 => y_in <= "10000011"; x_in <= "11001010"; z_correct<="0001101001011110";
        when 843 => y_in <= "10000011"; x_in <= "11001011"; z_correct<="0001100111100001";
        when 844 => y_in <= "10000011"; x_in <= "11001100"; z_correct<="0001100101100100";
        when 845 => y_in <= "10000011"; x_in <= "11001101"; z_correct<="0001100011100111";
        when 846 => y_in <= "10000011"; x_in <= "11001110"; z_correct<="0001100001101010";
        when 847 => y_in <= "10000011"; x_in <= "11001111"; z_correct<="0001011111101101";
        when 848 => y_in <= "10000011"; x_in <= "11010000"; z_correct<="0001011101110000";
        when 849 => y_in <= "10000011"; x_in <= "11010001"; z_correct<="0001011011110011";
        when 850 => y_in <= "10000011"; x_in <= "11010010"; z_correct<="0001011001110110";
        when 851 => y_in <= "10000011"; x_in <= "11010011"; z_correct<="0001010111111001";
        when 852 => y_in <= "10000011"; x_in <= "11010100"; z_correct<="0001010101111100";
        when 853 => y_in <= "10000011"; x_in <= "11010101"; z_correct<="0001010011111111";
        when 854 => y_in <= "10000011"; x_in <= "11010110"; z_correct<="0001010010000010";
        when 855 => y_in <= "10000011"; x_in <= "11010111"; z_correct<="0001010000000101";
        when 856 => y_in <= "10000011"; x_in <= "11011000"; z_correct<="0001001110001000";
        when 857 => y_in <= "10000011"; x_in <= "11011001"; z_correct<="0001001100001011";
        when 858 => y_in <= "10000011"; x_in <= "11011010"; z_correct<="0001001010001110";
        when 859 => y_in <= "10000011"; x_in <= "11011011"; z_correct<="0001001000010001";
        when 860 => y_in <= "10000011"; x_in <= "11011100"; z_correct<="0001000110010100";
        when 861 => y_in <= "10000011"; x_in <= "11011101"; z_correct<="0001000100010111";
        when 862 => y_in <= "10000011"; x_in <= "11011110"; z_correct<="0001000010011010";
        when 863 => y_in <= "10000011"; x_in <= "11011111"; z_correct<="0001000000011101";
        when 864 => y_in <= "10000011"; x_in <= "11100000"; z_correct<="0000111110100000";
        when 865 => y_in <= "10000011"; x_in <= "11100001"; z_correct<="0000111100100011";
        when 866 => y_in <= "10000011"; x_in <= "11100010"; z_correct<="0000111010100110";
        when 867 => y_in <= "10000011"; x_in <= "11100011"; z_correct<="0000111000101001";
        when 868 => y_in <= "10000011"; x_in <= "11100100"; z_correct<="0000110110101100";
        when 869 => y_in <= "10000011"; x_in <= "11100101"; z_correct<="0000110100101111";
        when 870 => y_in <= "10000011"; x_in <= "11100110"; z_correct<="0000110010110010";
        when 871 => y_in <= "10000011"; x_in <= "11100111"; z_correct<="0000110000110101";
        when 872 => y_in <= "10000011"; x_in <= "11101000"; z_correct<="0000101110111000";
        when 873 => y_in <= "10000011"; x_in <= "11101001"; z_correct<="0000101100111011";
        when 874 => y_in <= "10000011"; x_in <= "11101010"; z_correct<="0000101010111110";
        when 875 => y_in <= "10000011"; x_in <= "11101011"; z_correct<="0000101001000001";
        when 876 => y_in <= "10000011"; x_in <= "11101100"; z_correct<="0000100111000100";
        when 877 => y_in <= "10000011"; x_in <= "11101101"; z_correct<="0000100101000111";
        when 878 => y_in <= "10000011"; x_in <= "11101110"; z_correct<="0000100011001010";
        when 879 => y_in <= "10000011"; x_in <= "11101111"; z_correct<="0000100001001101";
        when 880 => y_in <= "10000011"; x_in <= "11110000"; z_correct<="0000011111010000";
        when 881 => y_in <= "10000011"; x_in <= "11110001"; z_correct<="0000011101010011";
        when 882 => y_in <= "10000011"; x_in <= "11110010"; z_correct<="0000011011010110";
        when 883 => y_in <= "10000011"; x_in <= "11110011"; z_correct<="0000011001011001";
        when 884 => y_in <= "10000011"; x_in <= "11110100"; z_correct<="0000010111011100";
        when 885 => y_in <= "10000011"; x_in <= "11110101"; z_correct<="0000010101011111";
        when 886 => y_in <= "10000011"; x_in <= "11110110"; z_correct<="0000010011100010";
        when 887 => y_in <= "10000011"; x_in <= "11110111"; z_correct<="0000010001100101";
        when 888 => y_in <= "10000011"; x_in <= "11111000"; z_correct<="0000001111101000";
        when 889 => y_in <= "10000011"; x_in <= "11111001"; z_correct<="0000001101101011";
        when 890 => y_in <= "10000011"; x_in <= "11111010"; z_correct<="0000001011101110";
        when 891 => y_in <= "10000011"; x_in <= "11111011"; z_correct<="0000001001110001";
        when 892 => y_in <= "10000011"; x_in <= "11111100"; z_correct<="0000000111110100";
        when 893 => y_in <= "10000011"; x_in <= "11111101"; z_correct<="0000000101110111";
        when 894 => y_in <= "10000011"; x_in <= "11111110"; z_correct<="0000000011111010";
        when 895 => y_in <= "10000011"; x_in <= "11111111"; z_correct<="0000000001111101";
        when 896 => y_in <= "10000011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 897 => y_in <= "10000011"; x_in <= "00000001"; z_correct<="1111111110000011";
        when 898 => y_in <= "10000011"; x_in <= "00000010"; z_correct<="1111111100000110";
        when 899 => y_in <= "10000011"; x_in <= "00000011"; z_correct<="1111111010001001";
        when 900 => y_in <= "10000011"; x_in <= "00000100"; z_correct<="1111111000001100";
        when 901 => y_in <= "10000011"; x_in <= "00000101"; z_correct<="1111110110001111";
        when 902 => y_in <= "10000011"; x_in <= "00000110"; z_correct<="1111110100010010";
        when 903 => y_in <= "10000011"; x_in <= "00000111"; z_correct<="1111110010010101";
        when 904 => y_in <= "10000011"; x_in <= "00001000"; z_correct<="1111110000011000";
        when 905 => y_in <= "10000011"; x_in <= "00001001"; z_correct<="1111101110011011";
        when 906 => y_in <= "10000011"; x_in <= "00001010"; z_correct<="1111101100011110";
        when 907 => y_in <= "10000011"; x_in <= "00001011"; z_correct<="1111101010100001";
        when 908 => y_in <= "10000011"; x_in <= "00001100"; z_correct<="1111101000100100";
        when 909 => y_in <= "10000011"; x_in <= "00001101"; z_correct<="1111100110100111";
        when 910 => y_in <= "10000011"; x_in <= "00001110"; z_correct<="1111100100101010";
        when 911 => y_in <= "10000011"; x_in <= "00001111"; z_correct<="1111100010101101";
        when 912 => y_in <= "10000011"; x_in <= "00010000"; z_correct<="1111100000110000";
        when 913 => y_in <= "10000011"; x_in <= "00010001"; z_correct<="1111011110110011";
        when 914 => y_in <= "10000011"; x_in <= "00010010"; z_correct<="1111011100110110";
        when 915 => y_in <= "10000011"; x_in <= "00010011"; z_correct<="1111011010111001";
        when 916 => y_in <= "10000011"; x_in <= "00010100"; z_correct<="1111011000111100";
        when 917 => y_in <= "10000011"; x_in <= "00010101"; z_correct<="1111010110111111";
        when 918 => y_in <= "10000011"; x_in <= "00010110"; z_correct<="1111010101000010";
        when 919 => y_in <= "10000011"; x_in <= "00010111"; z_correct<="1111010011000101";
        when 920 => y_in <= "10000011"; x_in <= "00011000"; z_correct<="1111010001001000";
        when 921 => y_in <= "10000011"; x_in <= "00011001"; z_correct<="1111001111001011";
        when 922 => y_in <= "10000011"; x_in <= "00011010"; z_correct<="1111001101001110";
        when 923 => y_in <= "10000011"; x_in <= "00011011"; z_correct<="1111001011010001";
        when 924 => y_in <= "10000011"; x_in <= "00011100"; z_correct<="1111001001010100";
        when 925 => y_in <= "10000011"; x_in <= "00011101"; z_correct<="1111000111010111";
        when 926 => y_in <= "10000011"; x_in <= "00011110"; z_correct<="1111000101011010";
        when 927 => y_in <= "10000011"; x_in <= "00011111"; z_correct<="1111000011011101";
        when 928 => y_in <= "10000011"; x_in <= "00100000"; z_correct<="1111000001100000";
        when 929 => y_in <= "10000011"; x_in <= "00100001"; z_correct<="1110111111100011";
        when 930 => y_in <= "10000011"; x_in <= "00100010"; z_correct<="1110111101100110";
        when 931 => y_in <= "10000011"; x_in <= "00100011"; z_correct<="1110111011101001";
        when 932 => y_in <= "10000011"; x_in <= "00100100"; z_correct<="1110111001101100";
        when 933 => y_in <= "10000011"; x_in <= "00100101"; z_correct<="1110110111101111";
        when 934 => y_in <= "10000011"; x_in <= "00100110"; z_correct<="1110110101110010";
        when 935 => y_in <= "10000011"; x_in <= "00100111"; z_correct<="1110110011110101";
        when 936 => y_in <= "10000011"; x_in <= "00101000"; z_correct<="1110110001111000";
        when 937 => y_in <= "10000011"; x_in <= "00101001"; z_correct<="1110101111111011";
        when 938 => y_in <= "10000011"; x_in <= "00101010"; z_correct<="1110101101111110";
        when 939 => y_in <= "10000011"; x_in <= "00101011"; z_correct<="1110101100000001";
        when 940 => y_in <= "10000011"; x_in <= "00101100"; z_correct<="1110101010000100";
        when 941 => y_in <= "10000011"; x_in <= "00101101"; z_correct<="1110101000000111";
        when 942 => y_in <= "10000011"; x_in <= "00101110"; z_correct<="1110100110001010";
        when 943 => y_in <= "10000011"; x_in <= "00101111"; z_correct<="1110100100001101";
        when 944 => y_in <= "10000011"; x_in <= "00110000"; z_correct<="1110100010010000";
        when 945 => y_in <= "10000011"; x_in <= "00110001"; z_correct<="1110100000010011";
        when 946 => y_in <= "10000011"; x_in <= "00110010"; z_correct<="1110011110010110";
        when 947 => y_in <= "10000011"; x_in <= "00110011"; z_correct<="1110011100011001";
        when 948 => y_in <= "10000011"; x_in <= "00110100"; z_correct<="1110011010011100";
        when 949 => y_in <= "10000011"; x_in <= "00110101"; z_correct<="1110011000011111";
        when 950 => y_in <= "10000011"; x_in <= "00110110"; z_correct<="1110010110100010";
        when 951 => y_in <= "10000011"; x_in <= "00110111"; z_correct<="1110010100100101";
        when 952 => y_in <= "10000011"; x_in <= "00111000"; z_correct<="1110010010101000";
        when 953 => y_in <= "10000011"; x_in <= "00111001"; z_correct<="1110010000101011";
        when 954 => y_in <= "10000011"; x_in <= "00111010"; z_correct<="1110001110101110";
        when 955 => y_in <= "10000011"; x_in <= "00111011"; z_correct<="1110001100110001";
        when 956 => y_in <= "10000011"; x_in <= "00111100"; z_correct<="1110001010110100";
        when 957 => y_in <= "10000011"; x_in <= "00111101"; z_correct<="1110001000110111";
        when 958 => y_in <= "10000011"; x_in <= "00111110"; z_correct<="1110000110111010";
        when 959 => y_in <= "10000011"; x_in <= "00111111"; z_correct<="1110000100111101";
        when 960 => y_in <= "10000011"; x_in <= "01000000"; z_correct<="1110000011000000";
        when 961 => y_in <= "10000011"; x_in <= "01000001"; z_correct<="1110000001000011";
        when 962 => y_in <= "10000011"; x_in <= "01000010"; z_correct<="1101111111000110";
        when 963 => y_in <= "10000011"; x_in <= "01000011"; z_correct<="1101111101001001";
        when 964 => y_in <= "10000011"; x_in <= "01000100"; z_correct<="1101111011001100";
        when 965 => y_in <= "10000011"; x_in <= "01000101"; z_correct<="1101111001001111";
        when 966 => y_in <= "10000011"; x_in <= "01000110"; z_correct<="1101110111010010";
        when 967 => y_in <= "10000011"; x_in <= "01000111"; z_correct<="1101110101010101";
        when 968 => y_in <= "10000011"; x_in <= "01001000"; z_correct<="1101110011011000";
        when 969 => y_in <= "10000011"; x_in <= "01001001"; z_correct<="1101110001011011";
        when 970 => y_in <= "10000011"; x_in <= "01001010"; z_correct<="1101101111011110";
        when 971 => y_in <= "10000011"; x_in <= "01001011"; z_correct<="1101101101100001";
        when 972 => y_in <= "10000011"; x_in <= "01001100"; z_correct<="1101101011100100";
        when 973 => y_in <= "10000011"; x_in <= "01001101"; z_correct<="1101101001100111";
        when 974 => y_in <= "10000011"; x_in <= "01001110"; z_correct<="1101100111101010";
        when 975 => y_in <= "10000011"; x_in <= "01001111"; z_correct<="1101100101101101";
        when 976 => y_in <= "10000011"; x_in <= "01010000"; z_correct<="1101100011110000";
        when 977 => y_in <= "10000011"; x_in <= "01010001"; z_correct<="1101100001110011";
        when 978 => y_in <= "10000011"; x_in <= "01010010"; z_correct<="1101011111110110";
        when 979 => y_in <= "10000011"; x_in <= "01010011"; z_correct<="1101011101111001";
        when 980 => y_in <= "10000011"; x_in <= "01010100"; z_correct<="1101011011111100";
        when 981 => y_in <= "10000011"; x_in <= "01010101"; z_correct<="1101011001111111";
        when 982 => y_in <= "10000011"; x_in <= "01010110"; z_correct<="1101011000000010";
        when 983 => y_in <= "10000011"; x_in <= "01010111"; z_correct<="1101010110000101";
        when 984 => y_in <= "10000011"; x_in <= "01011000"; z_correct<="1101010100001000";
        when 985 => y_in <= "10000011"; x_in <= "01011001"; z_correct<="1101010010001011";
        when 986 => y_in <= "10000011"; x_in <= "01011010"; z_correct<="1101010000001110";
        when 987 => y_in <= "10000011"; x_in <= "01011011"; z_correct<="1101001110010001";
        when 988 => y_in <= "10000011"; x_in <= "01011100"; z_correct<="1101001100010100";
        when 989 => y_in <= "10000011"; x_in <= "01011101"; z_correct<="1101001010010111";
        when 990 => y_in <= "10000011"; x_in <= "01011110"; z_correct<="1101001000011010";
        when 991 => y_in <= "10000011"; x_in <= "01011111"; z_correct<="1101000110011101";
        when 992 => y_in <= "10000011"; x_in <= "01100000"; z_correct<="1101000100100000";
        when 993 => y_in <= "10000011"; x_in <= "01100001"; z_correct<="1101000010100011";
        when 994 => y_in <= "10000011"; x_in <= "01100010"; z_correct<="1101000000100110";
        when 995 => y_in <= "10000011"; x_in <= "01100011"; z_correct<="1100111110101001";
        when 996 => y_in <= "10000011"; x_in <= "01100100"; z_correct<="1100111100101100";
        when 997 => y_in <= "10000011"; x_in <= "01100101"; z_correct<="1100111010101111";
        when 998 => y_in <= "10000011"; x_in <= "01100110"; z_correct<="1100111000110010";
        when 999 => y_in <= "10000011"; x_in <= "01100111"; z_correct<="1100110110110101";
        when 1000 => y_in <= "10000011"; x_in <= "01101000"; z_correct<="1100110100111000";
        when 1001 => y_in <= "10000011"; x_in <= "01101001"; z_correct<="1100110010111011";
        when 1002 => y_in <= "10000011"; x_in <= "01101010"; z_correct<="1100110000111110";
        when 1003 => y_in <= "10000011"; x_in <= "01101011"; z_correct<="1100101111000001";
        when 1004 => y_in <= "10000011"; x_in <= "01101100"; z_correct<="1100101101000100";
        when 1005 => y_in <= "10000011"; x_in <= "01101101"; z_correct<="1100101011000111";
        when 1006 => y_in <= "10000011"; x_in <= "01101110"; z_correct<="1100101001001010";
        when 1007 => y_in <= "10000011"; x_in <= "01101111"; z_correct<="1100100111001101";
        when 1008 => y_in <= "10000011"; x_in <= "01110000"; z_correct<="1100100101010000";
        when 1009 => y_in <= "10000011"; x_in <= "01110001"; z_correct<="1100100011010011";
        when 1010 => y_in <= "10000011"; x_in <= "01110010"; z_correct<="1100100001010110";
        when 1011 => y_in <= "10000011"; x_in <= "01110011"; z_correct<="1100011111011001";
        when 1012 => y_in <= "10000011"; x_in <= "01110100"; z_correct<="1100011101011100";
        when 1013 => y_in <= "10000011"; x_in <= "01110101"; z_correct<="1100011011011111";
        when 1014 => y_in <= "10000011"; x_in <= "01110110"; z_correct<="1100011001100010";
        when 1015 => y_in <= "10000011"; x_in <= "01110111"; z_correct<="1100010111100101";
        when 1016 => y_in <= "10000011"; x_in <= "01111000"; z_correct<="1100010101101000";
        when 1017 => y_in <= "10000011"; x_in <= "01111001"; z_correct<="1100010011101011";
        when 1018 => y_in <= "10000011"; x_in <= "01111010"; z_correct<="1100010001101110";
        when 1019 => y_in <= "10000011"; x_in <= "01111011"; z_correct<="1100001111110001";
        when 1020 => y_in <= "10000011"; x_in <= "01111100"; z_correct<="1100001101110100";
        when 1021 => y_in <= "10000011"; x_in <= "01111101"; z_correct<="1100001011110111";
        when 1022 => y_in <= "10000011"; x_in <= "01111110"; z_correct<="1100001001111010";
        when 1023 => y_in <= "10000011"; x_in <= "01111111"; z_correct<="1100000111111101";
        when 1024 => y_in <= "10000100"; x_in <= "10000000"; z_correct<="0011111000000000";
        when 1025 => y_in <= "10000100"; x_in <= "10000001"; z_correct<="0011110110000100";
        when 1026 => y_in <= "10000100"; x_in <= "10000010"; z_correct<="0011110100001000";
        when 1027 => y_in <= "10000100"; x_in <= "10000011"; z_correct<="0011110010001100";
        when 1028 => y_in <= "10000100"; x_in <= "10000100"; z_correct<="0011110000010000";
        when 1029 => y_in <= "10000100"; x_in <= "10000101"; z_correct<="0011101110010100";
        when 1030 => y_in <= "10000100"; x_in <= "10000110"; z_correct<="0011101100011000";
        when 1031 => y_in <= "10000100"; x_in <= "10000111"; z_correct<="0011101010011100";
        when 1032 => y_in <= "10000100"; x_in <= "10001000"; z_correct<="0011101000100000";
        when 1033 => y_in <= "10000100"; x_in <= "10001001"; z_correct<="0011100110100100";
        when 1034 => y_in <= "10000100"; x_in <= "10001010"; z_correct<="0011100100101000";
        when 1035 => y_in <= "10000100"; x_in <= "10001011"; z_correct<="0011100010101100";
        when 1036 => y_in <= "10000100"; x_in <= "10001100"; z_correct<="0011100000110000";
        when 1037 => y_in <= "10000100"; x_in <= "10001101"; z_correct<="0011011110110100";
        when 1038 => y_in <= "10000100"; x_in <= "10001110"; z_correct<="0011011100111000";
        when 1039 => y_in <= "10000100"; x_in <= "10001111"; z_correct<="0011011010111100";
        when 1040 => y_in <= "10000100"; x_in <= "10010000"; z_correct<="0011011001000000";
        when 1041 => y_in <= "10000100"; x_in <= "10010001"; z_correct<="0011010111000100";
        when 1042 => y_in <= "10000100"; x_in <= "10010010"; z_correct<="0011010101001000";
        when 1043 => y_in <= "10000100"; x_in <= "10010011"; z_correct<="0011010011001100";
        when 1044 => y_in <= "10000100"; x_in <= "10010100"; z_correct<="0011010001010000";
        when 1045 => y_in <= "10000100"; x_in <= "10010101"; z_correct<="0011001111010100";
        when 1046 => y_in <= "10000100"; x_in <= "10010110"; z_correct<="0011001101011000";
        when 1047 => y_in <= "10000100"; x_in <= "10010111"; z_correct<="0011001011011100";
        when 1048 => y_in <= "10000100"; x_in <= "10011000"; z_correct<="0011001001100000";
        when 1049 => y_in <= "10000100"; x_in <= "10011001"; z_correct<="0011000111100100";
        when 1050 => y_in <= "10000100"; x_in <= "10011010"; z_correct<="0011000101101000";
        when 1051 => y_in <= "10000100"; x_in <= "10011011"; z_correct<="0011000011101100";
        when 1052 => y_in <= "10000100"; x_in <= "10011100"; z_correct<="0011000001110000";
        when 1053 => y_in <= "10000100"; x_in <= "10011101"; z_correct<="0010111111110100";
        when 1054 => y_in <= "10000100"; x_in <= "10011110"; z_correct<="0010111101111000";
        when 1055 => y_in <= "10000100"; x_in <= "10011111"; z_correct<="0010111011111100";
        when 1056 => y_in <= "10000100"; x_in <= "10100000"; z_correct<="0010111010000000";
        when 1057 => y_in <= "10000100"; x_in <= "10100001"; z_correct<="0010111000000100";
        when 1058 => y_in <= "10000100"; x_in <= "10100010"; z_correct<="0010110110001000";
        when 1059 => y_in <= "10000100"; x_in <= "10100011"; z_correct<="0010110100001100";
        when 1060 => y_in <= "10000100"; x_in <= "10100100"; z_correct<="0010110010010000";
        when 1061 => y_in <= "10000100"; x_in <= "10100101"; z_correct<="0010110000010100";
        when 1062 => y_in <= "10000100"; x_in <= "10100110"; z_correct<="0010101110011000";
        when 1063 => y_in <= "10000100"; x_in <= "10100111"; z_correct<="0010101100011100";
        when 1064 => y_in <= "10000100"; x_in <= "10101000"; z_correct<="0010101010100000";
        when 1065 => y_in <= "10000100"; x_in <= "10101001"; z_correct<="0010101000100100";
        when 1066 => y_in <= "10000100"; x_in <= "10101010"; z_correct<="0010100110101000";
        when 1067 => y_in <= "10000100"; x_in <= "10101011"; z_correct<="0010100100101100";
        when 1068 => y_in <= "10000100"; x_in <= "10101100"; z_correct<="0010100010110000";
        when 1069 => y_in <= "10000100"; x_in <= "10101101"; z_correct<="0010100000110100";
        when 1070 => y_in <= "10000100"; x_in <= "10101110"; z_correct<="0010011110111000";
        when 1071 => y_in <= "10000100"; x_in <= "10101111"; z_correct<="0010011100111100";
        when 1072 => y_in <= "10000100"; x_in <= "10110000"; z_correct<="0010011011000000";
        when 1073 => y_in <= "10000100"; x_in <= "10110001"; z_correct<="0010011001000100";
        when 1074 => y_in <= "10000100"; x_in <= "10110010"; z_correct<="0010010111001000";
        when 1075 => y_in <= "10000100"; x_in <= "10110011"; z_correct<="0010010101001100";
        when 1076 => y_in <= "10000100"; x_in <= "10110100"; z_correct<="0010010011010000";
        when 1077 => y_in <= "10000100"; x_in <= "10110101"; z_correct<="0010010001010100";
        when 1078 => y_in <= "10000100"; x_in <= "10110110"; z_correct<="0010001111011000";
        when 1079 => y_in <= "10000100"; x_in <= "10110111"; z_correct<="0010001101011100";
        when 1080 => y_in <= "10000100"; x_in <= "10111000"; z_correct<="0010001011100000";
        when 1081 => y_in <= "10000100"; x_in <= "10111001"; z_correct<="0010001001100100";
        when 1082 => y_in <= "10000100"; x_in <= "10111010"; z_correct<="0010000111101000";
        when 1083 => y_in <= "10000100"; x_in <= "10111011"; z_correct<="0010000101101100";
        when 1084 => y_in <= "10000100"; x_in <= "10111100"; z_correct<="0010000011110000";
        when 1085 => y_in <= "10000100"; x_in <= "10111101"; z_correct<="0010000001110100";
        when 1086 => y_in <= "10000100"; x_in <= "10111110"; z_correct<="0001111111111000";
        when 1087 => y_in <= "10000100"; x_in <= "10111111"; z_correct<="0001111101111100";
        when 1088 => y_in <= "10000100"; x_in <= "11000000"; z_correct<="0001111100000000";
        when 1089 => y_in <= "10000100"; x_in <= "11000001"; z_correct<="0001111010000100";
        when 1090 => y_in <= "10000100"; x_in <= "11000010"; z_correct<="0001111000001000";
        when 1091 => y_in <= "10000100"; x_in <= "11000011"; z_correct<="0001110110001100";
        when 1092 => y_in <= "10000100"; x_in <= "11000100"; z_correct<="0001110100010000";
        when 1093 => y_in <= "10000100"; x_in <= "11000101"; z_correct<="0001110010010100";
        when 1094 => y_in <= "10000100"; x_in <= "11000110"; z_correct<="0001110000011000";
        when 1095 => y_in <= "10000100"; x_in <= "11000111"; z_correct<="0001101110011100";
        when 1096 => y_in <= "10000100"; x_in <= "11001000"; z_correct<="0001101100100000";
        when 1097 => y_in <= "10000100"; x_in <= "11001001"; z_correct<="0001101010100100";
        when 1098 => y_in <= "10000100"; x_in <= "11001010"; z_correct<="0001101000101000";
        when 1099 => y_in <= "10000100"; x_in <= "11001011"; z_correct<="0001100110101100";
        when 1100 => y_in <= "10000100"; x_in <= "11001100"; z_correct<="0001100100110000";
        when 1101 => y_in <= "10000100"; x_in <= "11001101"; z_correct<="0001100010110100";
        when 1102 => y_in <= "10000100"; x_in <= "11001110"; z_correct<="0001100000111000";
        when 1103 => y_in <= "10000100"; x_in <= "11001111"; z_correct<="0001011110111100";
        when 1104 => y_in <= "10000100"; x_in <= "11010000"; z_correct<="0001011101000000";
        when 1105 => y_in <= "10000100"; x_in <= "11010001"; z_correct<="0001011011000100";
        when 1106 => y_in <= "10000100"; x_in <= "11010010"; z_correct<="0001011001001000";
        when 1107 => y_in <= "10000100"; x_in <= "11010011"; z_correct<="0001010111001100";
        when 1108 => y_in <= "10000100"; x_in <= "11010100"; z_correct<="0001010101010000";
        when 1109 => y_in <= "10000100"; x_in <= "11010101"; z_correct<="0001010011010100";
        when 1110 => y_in <= "10000100"; x_in <= "11010110"; z_correct<="0001010001011000";
        when 1111 => y_in <= "10000100"; x_in <= "11010111"; z_correct<="0001001111011100";
        when 1112 => y_in <= "10000100"; x_in <= "11011000"; z_correct<="0001001101100000";
        when 1113 => y_in <= "10000100"; x_in <= "11011001"; z_correct<="0001001011100100";
        when 1114 => y_in <= "10000100"; x_in <= "11011010"; z_correct<="0001001001101000";
        when 1115 => y_in <= "10000100"; x_in <= "11011011"; z_correct<="0001000111101100";
        when 1116 => y_in <= "10000100"; x_in <= "11011100"; z_correct<="0001000101110000";
        when 1117 => y_in <= "10000100"; x_in <= "11011101"; z_correct<="0001000011110100";
        when 1118 => y_in <= "10000100"; x_in <= "11011110"; z_correct<="0001000001111000";
        when 1119 => y_in <= "10000100"; x_in <= "11011111"; z_correct<="0000111111111100";
        when 1120 => y_in <= "10000100"; x_in <= "11100000"; z_correct<="0000111110000000";
        when 1121 => y_in <= "10000100"; x_in <= "11100001"; z_correct<="0000111100000100";
        when 1122 => y_in <= "10000100"; x_in <= "11100010"; z_correct<="0000111010001000";
        when 1123 => y_in <= "10000100"; x_in <= "11100011"; z_correct<="0000111000001100";
        when 1124 => y_in <= "10000100"; x_in <= "11100100"; z_correct<="0000110110010000";
        when 1125 => y_in <= "10000100"; x_in <= "11100101"; z_correct<="0000110100010100";
        when 1126 => y_in <= "10000100"; x_in <= "11100110"; z_correct<="0000110010011000";
        when 1127 => y_in <= "10000100"; x_in <= "11100111"; z_correct<="0000110000011100";
        when 1128 => y_in <= "10000100"; x_in <= "11101000"; z_correct<="0000101110100000";
        when 1129 => y_in <= "10000100"; x_in <= "11101001"; z_correct<="0000101100100100";
        when 1130 => y_in <= "10000100"; x_in <= "11101010"; z_correct<="0000101010101000";
        when 1131 => y_in <= "10000100"; x_in <= "11101011"; z_correct<="0000101000101100";
        when 1132 => y_in <= "10000100"; x_in <= "11101100"; z_correct<="0000100110110000";
        when 1133 => y_in <= "10000100"; x_in <= "11101101"; z_correct<="0000100100110100";
        when 1134 => y_in <= "10000100"; x_in <= "11101110"; z_correct<="0000100010111000";
        when 1135 => y_in <= "10000100"; x_in <= "11101111"; z_correct<="0000100000111100";
        when 1136 => y_in <= "10000100"; x_in <= "11110000"; z_correct<="0000011111000000";
        when 1137 => y_in <= "10000100"; x_in <= "11110001"; z_correct<="0000011101000100";
        when 1138 => y_in <= "10000100"; x_in <= "11110010"; z_correct<="0000011011001000";
        when 1139 => y_in <= "10000100"; x_in <= "11110011"; z_correct<="0000011001001100";
        when 1140 => y_in <= "10000100"; x_in <= "11110100"; z_correct<="0000010111010000";
        when 1141 => y_in <= "10000100"; x_in <= "11110101"; z_correct<="0000010101010100";
        when 1142 => y_in <= "10000100"; x_in <= "11110110"; z_correct<="0000010011011000";
        when 1143 => y_in <= "10000100"; x_in <= "11110111"; z_correct<="0000010001011100";
        when 1144 => y_in <= "10000100"; x_in <= "11111000"; z_correct<="0000001111100000";
        when 1145 => y_in <= "10000100"; x_in <= "11111001"; z_correct<="0000001101100100";
        when 1146 => y_in <= "10000100"; x_in <= "11111010"; z_correct<="0000001011101000";
        when 1147 => y_in <= "10000100"; x_in <= "11111011"; z_correct<="0000001001101100";
        when 1148 => y_in <= "10000100"; x_in <= "11111100"; z_correct<="0000000111110000";
        when 1149 => y_in <= "10000100"; x_in <= "11111101"; z_correct<="0000000101110100";
        when 1150 => y_in <= "10000100"; x_in <= "11111110"; z_correct<="0000000011111000";
        when 1151 => y_in <= "10000100"; x_in <= "11111111"; z_correct<="0000000001111100";
        when 1152 => y_in <= "10000100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 1153 => y_in <= "10000100"; x_in <= "00000001"; z_correct<="1111111110000100";
        when 1154 => y_in <= "10000100"; x_in <= "00000010"; z_correct<="1111111100001000";
        when 1155 => y_in <= "10000100"; x_in <= "00000011"; z_correct<="1111111010001100";
        when 1156 => y_in <= "10000100"; x_in <= "00000100"; z_correct<="1111111000010000";
        when 1157 => y_in <= "10000100"; x_in <= "00000101"; z_correct<="1111110110010100";
        when 1158 => y_in <= "10000100"; x_in <= "00000110"; z_correct<="1111110100011000";
        when 1159 => y_in <= "10000100"; x_in <= "00000111"; z_correct<="1111110010011100";
        when 1160 => y_in <= "10000100"; x_in <= "00001000"; z_correct<="1111110000100000";
        when 1161 => y_in <= "10000100"; x_in <= "00001001"; z_correct<="1111101110100100";
        when 1162 => y_in <= "10000100"; x_in <= "00001010"; z_correct<="1111101100101000";
        when 1163 => y_in <= "10000100"; x_in <= "00001011"; z_correct<="1111101010101100";
        when 1164 => y_in <= "10000100"; x_in <= "00001100"; z_correct<="1111101000110000";
        when 1165 => y_in <= "10000100"; x_in <= "00001101"; z_correct<="1111100110110100";
        when 1166 => y_in <= "10000100"; x_in <= "00001110"; z_correct<="1111100100111000";
        when 1167 => y_in <= "10000100"; x_in <= "00001111"; z_correct<="1111100010111100";
        when 1168 => y_in <= "10000100"; x_in <= "00010000"; z_correct<="1111100001000000";
        when 1169 => y_in <= "10000100"; x_in <= "00010001"; z_correct<="1111011111000100";
        when 1170 => y_in <= "10000100"; x_in <= "00010010"; z_correct<="1111011101001000";
        when 1171 => y_in <= "10000100"; x_in <= "00010011"; z_correct<="1111011011001100";
        when 1172 => y_in <= "10000100"; x_in <= "00010100"; z_correct<="1111011001010000";
        when 1173 => y_in <= "10000100"; x_in <= "00010101"; z_correct<="1111010111010100";
        when 1174 => y_in <= "10000100"; x_in <= "00010110"; z_correct<="1111010101011000";
        when 1175 => y_in <= "10000100"; x_in <= "00010111"; z_correct<="1111010011011100";
        when 1176 => y_in <= "10000100"; x_in <= "00011000"; z_correct<="1111010001100000";
        when 1177 => y_in <= "10000100"; x_in <= "00011001"; z_correct<="1111001111100100";
        when 1178 => y_in <= "10000100"; x_in <= "00011010"; z_correct<="1111001101101000";
        when 1179 => y_in <= "10000100"; x_in <= "00011011"; z_correct<="1111001011101100";
        when 1180 => y_in <= "10000100"; x_in <= "00011100"; z_correct<="1111001001110000";
        when 1181 => y_in <= "10000100"; x_in <= "00011101"; z_correct<="1111000111110100";
        when 1182 => y_in <= "10000100"; x_in <= "00011110"; z_correct<="1111000101111000";
        when 1183 => y_in <= "10000100"; x_in <= "00011111"; z_correct<="1111000011111100";
        when 1184 => y_in <= "10000100"; x_in <= "00100000"; z_correct<="1111000010000000";
        when 1185 => y_in <= "10000100"; x_in <= "00100001"; z_correct<="1111000000000100";
        when 1186 => y_in <= "10000100"; x_in <= "00100010"; z_correct<="1110111110001000";
        when 1187 => y_in <= "10000100"; x_in <= "00100011"; z_correct<="1110111100001100";
        when 1188 => y_in <= "10000100"; x_in <= "00100100"; z_correct<="1110111010010000";
        when 1189 => y_in <= "10000100"; x_in <= "00100101"; z_correct<="1110111000010100";
        when 1190 => y_in <= "10000100"; x_in <= "00100110"; z_correct<="1110110110011000";
        when 1191 => y_in <= "10000100"; x_in <= "00100111"; z_correct<="1110110100011100";
        when 1192 => y_in <= "10000100"; x_in <= "00101000"; z_correct<="1110110010100000";
        when 1193 => y_in <= "10000100"; x_in <= "00101001"; z_correct<="1110110000100100";
        when 1194 => y_in <= "10000100"; x_in <= "00101010"; z_correct<="1110101110101000";
        when 1195 => y_in <= "10000100"; x_in <= "00101011"; z_correct<="1110101100101100";
        when 1196 => y_in <= "10000100"; x_in <= "00101100"; z_correct<="1110101010110000";
        when 1197 => y_in <= "10000100"; x_in <= "00101101"; z_correct<="1110101000110100";
        when 1198 => y_in <= "10000100"; x_in <= "00101110"; z_correct<="1110100110111000";
        when 1199 => y_in <= "10000100"; x_in <= "00101111"; z_correct<="1110100100111100";
        when 1200 => y_in <= "10000100"; x_in <= "00110000"; z_correct<="1110100011000000";
        when 1201 => y_in <= "10000100"; x_in <= "00110001"; z_correct<="1110100001000100";
        when 1202 => y_in <= "10000100"; x_in <= "00110010"; z_correct<="1110011111001000";
        when 1203 => y_in <= "10000100"; x_in <= "00110011"; z_correct<="1110011101001100";
        when 1204 => y_in <= "10000100"; x_in <= "00110100"; z_correct<="1110011011010000";
        when 1205 => y_in <= "10000100"; x_in <= "00110101"; z_correct<="1110011001010100";
        when 1206 => y_in <= "10000100"; x_in <= "00110110"; z_correct<="1110010111011000";
        when 1207 => y_in <= "10000100"; x_in <= "00110111"; z_correct<="1110010101011100";
        when 1208 => y_in <= "10000100"; x_in <= "00111000"; z_correct<="1110010011100000";
        when 1209 => y_in <= "10000100"; x_in <= "00111001"; z_correct<="1110010001100100";
        when 1210 => y_in <= "10000100"; x_in <= "00111010"; z_correct<="1110001111101000";
        when 1211 => y_in <= "10000100"; x_in <= "00111011"; z_correct<="1110001101101100";
        when 1212 => y_in <= "10000100"; x_in <= "00111100"; z_correct<="1110001011110000";
        when 1213 => y_in <= "10000100"; x_in <= "00111101"; z_correct<="1110001001110100";
        when 1214 => y_in <= "10000100"; x_in <= "00111110"; z_correct<="1110000111111000";
        when 1215 => y_in <= "10000100"; x_in <= "00111111"; z_correct<="1110000101111100";
        when 1216 => y_in <= "10000100"; x_in <= "01000000"; z_correct<="1110000100000000";
        when 1217 => y_in <= "10000100"; x_in <= "01000001"; z_correct<="1110000010000100";
        when 1218 => y_in <= "10000100"; x_in <= "01000010"; z_correct<="1110000000001000";
        when 1219 => y_in <= "10000100"; x_in <= "01000011"; z_correct<="1101111110001100";
        when 1220 => y_in <= "10000100"; x_in <= "01000100"; z_correct<="1101111100010000";
        when 1221 => y_in <= "10000100"; x_in <= "01000101"; z_correct<="1101111010010100";
        when 1222 => y_in <= "10000100"; x_in <= "01000110"; z_correct<="1101111000011000";
        when 1223 => y_in <= "10000100"; x_in <= "01000111"; z_correct<="1101110110011100";
        when 1224 => y_in <= "10000100"; x_in <= "01001000"; z_correct<="1101110100100000";
        when 1225 => y_in <= "10000100"; x_in <= "01001001"; z_correct<="1101110010100100";
        when 1226 => y_in <= "10000100"; x_in <= "01001010"; z_correct<="1101110000101000";
        when 1227 => y_in <= "10000100"; x_in <= "01001011"; z_correct<="1101101110101100";
        when 1228 => y_in <= "10000100"; x_in <= "01001100"; z_correct<="1101101100110000";
        when 1229 => y_in <= "10000100"; x_in <= "01001101"; z_correct<="1101101010110100";
        when 1230 => y_in <= "10000100"; x_in <= "01001110"; z_correct<="1101101000111000";
        when 1231 => y_in <= "10000100"; x_in <= "01001111"; z_correct<="1101100110111100";
        when 1232 => y_in <= "10000100"; x_in <= "01010000"; z_correct<="1101100101000000";
        when 1233 => y_in <= "10000100"; x_in <= "01010001"; z_correct<="1101100011000100";
        when 1234 => y_in <= "10000100"; x_in <= "01010010"; z_correct<="1101100001001000";
        when 1235 => y_in <= "10000100"; x_in <= "01010011"; z_correct<="1101011111001100";
        when 1236 => y_in <= "10000100"; x_in <= "01010100"; z_correct<="1101011101010000";
        when 1237 => y_in <= "10000100"; x_in <= "01010101"; z_correct<="1101011011010100";
        when 1238 => y_in <= "10000100"; x_in <= "01010110"; z_correct<="1101011001011000";
        when 1239 => y_in <= "10000100"; x_in <= "01010111"; z_correct<="1101010111011100";
        when 1240 => y_in <= "10000100"; x_in <= "01011000"; z_correct<="1101010101100000";
        when 1241 => y_in <= "10000100"; x_in <= "01011001"; z_correct<="1101010011100100";
        when 1242 => y_in <= "10000100"; x_in <= "01011010"; z_correct<="1101010001101000";
        when 1243 => y_in <= "10000100"; x_in <= "01011011"; z_correct<="1101001111101100";
        when 1244 => y_in <= "10000100"; x_in <= "01011100"; z_correct<="1101001101110000";
        when 1245 => y_in <= "10000100"; x_in <= "01011101"; z_correct<="1101001011110100";
        when 1246 => y_in <= "10000100"; x_in <= "01011110"; z_correct<="1101001001111000";
        when 1247 => y_in <= "10000100"; x_in <= "01011111"; z_correct<="1101000111111100";
        when 1248 => y_in <= "10000100"; x_in <= "01100000"; z_correct<="1101000110000000";
        when 1249 => y_in <= "10000100"; x_in <= "01100001"; z_correct<="1101000100000100";
        when 1250 => y_in <= "10000100"; x_in <= "01100010"; z_correct<="1101000010001000";
        when 1251 => y_in <= "10000100"; x_in <= "01100011"; z_correct<="1101000000001100";
        when 1252 => y_in <= "10000100"; x_in <= "01100100"; z_correct<="1100111110010000";
        when 1253 => y_in <= "10000100"; x_in <= "01100101"; z_correct<="1100111100010100";
        when 1254 => y_in <= "10000100"; x_in <= "01100110"; z_correct<="1100111010011000";
        when 1255 => y_in <= "10000100"; x_in <= "01100111"; z_correct<="1100111000011100";
        when 1256 => y_in <= "10000100"; x_in <= "01101000"; z_correct<="1100110110100000";
        when 1257 => y_in <= "10000100"; x_in <= "01101001"; z_correct<="1100110100100100";
        when 1258 => y_in <= "10000100"; x_in <= "01101010"; z_correct<="1100110010101000";
        when 1259 => y_in <= "10000100"; x_in <= "01101011"; z_correct<="1100110000101100";
        when 1260 => y_in <= "10000100"; x_in <= "01101100"; z_correct<="1100101110110000";
        when 1261 => y_in <= "10000100"; x_in <= "01101101"; z_correct<="1100101100110100";
        when 1262 => y_in <= "10000100"; x_in <= "01101110"; z_correct<="1100101010111000";
        when 1263 => y_in <= "10000100"; x_in <= "01101111"; z_correct<="1100101000111100";
        when 1264 => y_in <= "10000100"; x_in <= "01110000"; z_correct<="1100100111000000";
        when 1265 => y_in <= "10000100"; x_in <= "01110001"; z_correct<="1100100101000100";
        when 1266 => y_in <= "10000100"; x_in <= "01110010"; z_correct<="1100100011001000";
        when 1267 => y_in <= "10000100"; x_in <= "01110011"; z_correct<="1100100001001100";
        when 1268 => y_in <= "10000100"; x_in <= "01110100"; z_correct<="1100011111010000";
        when 1269 => y_in <= "10000100"; x_in <= "01110101"; z_correct<="1100011101010100";
        when 1270 => y_in <= "10000100"; x_in <= "01110110"; z_correct<="1100011011011000";
        when 1271 => y_in <= "10000100"; x_in <= "01110111"; z_correct<="1100011001011100";
        when 1272 => y_in <= "10000100"; x_in <= "01111000"; z_correct<="1100010111100000";
        when 1273 => y_in <= "10000100"; x_in <= "01111001"; z_correct<="1100010101100100";
        when 1274 => y_in <= "10000100"; x_in <= "01111010"; z_correct<="1100010011101000";
        when 1275 => y_in <= "10000100"; x_in <= "01111011"; z_correct<="1100010001101100";
        when 1276 => y_in <= "10000100"; x_in <= "01111100"; z_correct<="1100001111110000";
        when 1277 => y_in <= "10000100"; x_in <= "01111101"; z_correct<="1100001101110100";
        when 1278 => y_in <= "10000100"; x_in <= "01111110"; z_correct<="1100001011111000";
        when 1279 => y_in <= "10000100"; x_in <= "01111111"; z_correct<="1100001001111100";
        when 1280 => y_in <= "10000101"; x_in <= "10000000"; z_correct<="0011110110000000";
        when 1281 => y_in <= "10000101"; x_in <= "10000001"; z_correct<="0011110100000101";
        when 1282 => y_in <= "10000101"; x_in <= "10000010"; z_correct<="0011110010001010";
        when 1283 => y_in <= "10000101"; x_in <= "10000011"; z_correct<="0011110000001111";
        when 1284 => y_in <= "10000101"; x_in <= "10000100"; z_correct<="0011101110010100";
        when 1285 => y_in <= "10000101"; x_in <= "10000101"; z_correct<="0011101100011001";
        when 1286 => y_in <= "10000101"; x_in <= "10000110"; z_correct<="0011101010011110";
        when 1287 => y_in <= "10000101"; x_in <= "10000111"; z_correct<="0011101000100011";
        when 1288 => y_in <= "10000101"; x_in <= "10001000"; z_correct<="0011100110101000";
        when 1289 => y_in <= "10000101"; x_in <= "10001001"; z_correct<="0011100100101101";
        when 1290 => y_in <= "10000101"; x_in <= "10001010"; z_correct<="0011100010110010";
        when 1291 => y_in <= "10000101"; x_in <= "10001011"; z_correct<="0011100000110111";
        when 1292 => y_in <= "10000101"; x_in <= "10001100"; z_correct<="0011011110111100";
        when 1293 => y_in <= "10000101"; x_in <= "10001101"; z_correct<="0011011101000001";
        when 1294 => y_in <= "10000101"; x_in <= "10001110"; z_correct<="0011011011000110";
        when 1295 => y_in <= "10000101"; x_in <= "10001111"; z_correct<="0011011001001011";
        when 1296 => y_in <= "10000101"; x_in <= "10010000"; z_correct<="0011010111010000";
        when 1297 => y_in <= "10000101"; x_in <= "10010001"; z_correct<="0011010101010101";
        when 1298 => y_in <= "10000101"; x_in <= "10010010"; z_correct<="0011010011011010";
        when 1299 => y_in <= "10000101"; x_in <= "10010011"; z_correct<="0011010001011111";
        when 1300 => y_in <= "10000101"; x_in <= "10010100"; z_correct<="0011001111100100";
        when 1301 => y_in <= "10000101"; x_in <= "10010101"; z_correct<="0011001101101001";
        when 1302 => y_in <= "10000101"; x_in <= "10010110"; z_correct<="0011001011101110";
        when 1303 => y_in <= "10000101"; x_in <= "10010111"; z_correct<="0011001001110011";
        when 1304 => y_in <= "10000101"; x_in <= "10011000"; z_correct<="0011000111111000";
        when 1305 => y_in <= "10000101"; x_in <= "10011001"; z_correct<="0011000101111101";
        when 1306 => y_in <= "10000101"; x_in <= "10011010"; z_correct<="0011000100000010";
        when 1307 => y_in <= "10000101"; x_in <= "10011011"; z_correct<="0011000010000111";
        when 1308 => y_in <= "10000101"; x_in <= "10011100"; z_correct<="0011000000001100";
        when 1309 => y_in <= "10000101"; x_in <= "10011101"; z_correct<="0010111110010001";
        when 1310 => y_in <= "10000101"; x_in <= "10011110"; z_correct<="0010111100010110";
        when 1311 => y_in <= "10000101"; x_in <= "10011111"; z_correct<="0010111010011011";
        when 1312 => y_in <= "10000101"; x_in <= "10100000"; z_correct<="0010111000100000";
        when 1313 => y_in <= "10000101"; x_in <= "10100001"; z_correct<="0010110110100101";
        when 1314 => y_in <= "10000101"; x_in <= "10100010"; z_correct<="0010110100101010";
        when 1315 => y_in <= "10000101"; x_in <= "10100011"; z_correct<="0010110010101111";
        when 1316 => y_in <= "10000101"; x_in <= "10100100"; z_correct<="0010110000110100";
        when 1317 => y_in <= "10000101"; x_in <= "10100101"; z_correct<="0010101110111001";
        when 1318 => y_in <= "10000101"; x_in <= "10100110"; z_correct<="0010101100111110";
        when 1319 => y_in <= "10000101"; x_in <= "10100111"; z_correct<="0010101011000011";
        when 1320 => y_in <= "10000101"; x_in <= "10101000"; z_correct<="0010101001001000";
        when 1321 => y_in <= "10000101"; x_in <= "10101001"; z_correct<="0010100111001101";
        when 1322 => y_in <= "10000101"; x_in <= "10101010"; z_correct<="0010100101010010";
        when 1323 => y_in <= "10000101"; x_in <= "10101011"; z_correct<="0010100011010111";
        when 1324 => y_in <= "10000101"; x_in <= "10101100"; z_correct<="0010100001011100";
        when 1325 => y_in <= "10000101"; x_in <= "10101101"; z_correct<="0010011111100001";
        when 1326 => y_in <= "10000101"; x_in <= "10101110"; z_correct<="0010011101100110";
        when 1327 => y_in <= "10000101"; x_in <= "10101111"; z_correct<="0010011011101011";
        when 1328 => y_in <= "10000101"; x_in <= "10110000"; z_correct<="0010011001110000";
        when 1329 => y_in <= "10000101"; x_in <= "10110001"; z_correct<="0010010111110101";
        when 1330 => y_in <= "10000101"; x_in <= "10110010"; z_correct<="0010010101111010";
        when 1331 => y_in <= "10000101"; x_in <= "10110011"; z_correct<="0010010011111111";
        when 1332 => y_in <= "10000101"; x_in <= "10110100"; z_correct<="0010010010000100";
        when 1333 => y_in <= "10000101"; x_in <= "10110101"; z_correct<="0010010000001001";
        when 1334 => y_in <= "10000101"; x_in <= "10110110"; z_correct<="0010001110001110";
        when 1335 => y_in <= "10000101"; x_in <= "10110111"; z_correct<="0010001100010011";
        when 1336 => y_in <= "10000101"; x_in <= "10111000"; z_correct<="0010001010011000";
        when 1337 => y_in <= "10000101"; x_in <= "10111001"; z_correct<="0010001000011101";
        when 1338 => y_in <= "10000101"; x_in <= "10111010"; z_correct<="0010000110100010";
        when 1339 => y_in <= "10000101"; x_in <= "10111011"; z_correct<="0010000100100111";
        when 1340 => y_in <= "10000101"; x_in <= "10111100"; z_correct<="0010000010101100";
        when 1341 => y_in <= "10000101"; x_in <= "10111101"; z_correct<="0010000000110001";
        when 1342 => y_in <= "10000101"; x_in <= "10111110"; z_correct<="0001111110110110";
        when 1343 => y_in <= "10000101"; x_in <= "10111111"; z_correct<="0001111100111011";
        when 1344 => y_in <= "10000101"; x_in <= "11000000"; z_correct<="0001111011000000";
        when 1345 => y_in <= "10000101"; x_in <= "11000001"; z_correct<="0001111001000101";
        when 1346 => y_in <= "10000101"; x_in <= "11000010"; z_correct<="0001110111001010";
        when 1347 => y_in <= "10000101"; x_in <= "11000011"; z_correct<="0001110101001111";
        when 1348 => y_in <= "10000101"; x_in <= "11000100"; z_correct<="0001110011010100";
        when 1349 => y_in <= "10000101"; x_in <= "11000101"; z_correct<="0001110001011001";
        when 1350 => y_in <= "10000101"; x_in <= "11000110"; z_correct<="0001101111011110";
        when 1351 => y_in <= "10000101"; x_in <= "11000111"; z_correct<="0001101101100011";
        when 1352 => y_in <= "10000101"; x_in <= "11001000"; z_correct<="0001101011101000";
        when 1353 => y_in <= "10000101"; x_in <= "11001001"; z_correct<="0001101001101101";
        when 1354 => y_in <= "10000101"; x_in <= "11001010"; z_correct<="0001100111110010";
        when 1355 => y_in <= "10000101"; x_in <= "11001011"; z_correct<="0001100101110111";
        when 1356 => y_in <= "10000101"; x_in <= "11001100"; z_correct<="0001100011111100";
        when 1357 => y_in <= "10000101"; x_in <= "11001101"; z_correct<="0001100010000001";
        when 1358 => y_in <= "10000101"; x_in <= "11001110"; z_correct<="0001100000000110";
        when 1359 => y_in <= "10000101"; x_in <= "11001111"; z_correct<="0001011110001011";
        when 1360 => y_in <= "10000101"; x_in <= "11010000"; z_correct<="0001011100010000";
        when 1361 => y_in <= "10000101"; x_in <= "11010001"; z_correct<="0001011010010101";
        when 1362 => y_in <= "10000101"; x_in <= "11010010"; z_correct<="0001011000011010";
        when 1363 => y_in <= "10000101"; x_in <= "11010011"; z_correct<="0001010110011111";
        when 1364 => y_in <= "10000101"; x_in <= "11010100"; z_correct<="0001010100100100";
        when 1365 => y_in <= "10000101"; x_in <= "11010101"; z_correct<="0001010010101001";
        when 1366 => y_in <= "10000101"; x_in <= "11010110"; z_correct<="0001010000101110";
        when 1367 => y_in <= "10000101"; x_in <= "11010111"; z_correct<="0001001110110011";
        when 1368 => y_in <= "10000101"; x_in <= "11011000"; z_correct<="0001001100111000";
        when 1369 => y_in <= "10000101"; x_in <= "11011001"; z_correct<="0001001010111101";
        when 1370 => y_in <= "10000101"; x_in <= "11011010"; z_correct<="0001001001000010";
        when 1371 => y_in <= "10000101"; x_in <= "11011011"; z_correct<="0001000111000111";
        when 1372 => y_in <= "10000101"; x_in <= "11011100"; z_correct<="0001000101001100";
        when 1373 => y_in <= "10000101"; x_in <= "11011101"; z_correct<="0001000011010001";
        when 1374 => y_in <= "10000101"; x_in <= "11011110"; z_correct<="0001000001010110";
        when 1375 => y_in <= "10000101"; x_in <= "11011111"; z_correct<="0000111111011011";
        when 1376 => y_in <= "10000101"; x_in <= "11100000"; z_correct<="0000111101100000";
        when 1377 => y_in <= "10000101"; x_in <= "11100001"; z_correct<="0000111011100101";
        when 1378 => y_in <= "10000101"; x_in <= "11100010"; z_correct<="0000111001101010";
        when 1379 => y_in <= "10000101"; x_in <= "11100011"; z_correct<="0000110111101111";
        when 1380 => y_in <= "10000101"; x_in <= "11100100"; z_correct<="0000110101110100";
        when 1381 => y_in <= "10000101"; x_in <= "11100101"; z_correct<="0000110011111001";
        when 1382 => y_in <= "10000101"; x_in <= "11100110"; z_correct<="0000110001111110";
        when 1383 => y_in <= "10000101"; x_in <= "11100111"; z_correct<="0000110000000011";
        when 1384 => y_in <= "10000101"; x_in <= "11101000"; z_correct<="0000101110001000";
        when 1385 => y_in <= "10000101"; x_in <= "11101001"; z_correct<="0000101100001101";
        when 1386 => y_in <= "10000101"; x_in <= "11101010"; z_correct<="0000101010010010";
        when 1387 => y_in <= "10000101"; x_in <= "11101011"; z_correct<="0000101000010111";
        when 1388 => y_in <= "10000101"; x_in <= "11101100"; z_correct<="0000100110011100";
        when 1389 => y_in <= "10000101"; x_in <= "11101101"; z_correct<="0000100100100001";
        when 1390 => y_in <= "10000101"; x_in <= "11101110"; z_correct<="0000100010100110";
        when 1391 => y_in <= "10000101"; x_in <= "11101111"; z_correct<="0000100000101011";
        when 1392 => y_in <= "10000101"; x_in <= "11110000"; z_correct<="0000011110110000";
        when 1393 => y_in <= "10000101"; x_in <= "11110001"; z_correct<="0000011100110101";
        when 1394 => y_in <= "10000101"; x_in <= "11110010"; z_correct<="0000011010111010";
        when 1395 => y_in <= "10000101"; x_in <= "11110011"; z_correct<="0000011000111111";
        when 1396 => y_in <= "10000101"; x_in <= "11110100"; z_correct<="0000010111000100";
        when 1397 => y_in <= "10000101"; x_in <= "11110101"; z_correct<="0000010101001001";
        when 1398 => y_in <= "10000101"; x_in <= "11110110"; z_correct<="0000010011001110";
        when 1399 => y_in <= "10000101"; x_in <= "11110111"; z_correct<="0000010001010011";
        when 1400 => y_in <= "10000101"; x_in <= "11111000"; z_correct<="0000001111011000";
        when 1401 => y_in <= "10000101"; x_in <= "11111001"; z_correct<="0000001101011101";
        when 1402 => y_in <= "10000101"; x_in <= "11111010"; z_correct<="0000001011100010";
        when 1403 => y_in <= "10000101"; x_in <= "11111011"; z_correct<="0000001001100111";
        when 1404 => y_in <= "10000101"; x_in <= "11111100"; z_correct<="0000000111101100";
        when 1405 => y_in <= "10000101"; x_in <= "11111101"; z_correct<="0000000101110001";
        when 1406 => y_in <= "10000101"; x_in <= "11111110"; z_correct<="0000000011110110";
        when 1407 => y_in <= "10000101"; x_in <= "11111111"; z_correct<="0000000001111011";
        when 1408 => y_in <= "10000101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 1409 => y_in <= "10000101"; x_in <= "00000001"; z_correct<="1111111110000101";
        when 1410 => y_in <= "10000101"; x_in <= "00000010"; z_correct<="1111111100001010";
        when 1411 => y_in <= "10000101"; x_in <= "00000011"; z_correct<="1111111010001111";
        when 1412 => y_in <= "10000101"; x_in <= "00000100"; z_correct<="1111111000010100";
        when 1413 => y_in <= "10000101"; x_in <= "00000101"; z_correct<="1111110110011001";
        when 1414 => y_in <= "10000101"; x_in <= "00000110"; z_correct<="1111110100011110";
        when 1415 => y_in <= "10000101"; x_in <= "00000111"; z_correct<="1111110010100011";
        when 1416 => y_in <= "10000101"; x_in <= "00001000"; z_correct<="1111110000101000";
        when 1417 => y_in <= "10000101"; x_in <= "00001001"; z_correct<="1111101110101101";
        when 1418 => y_in <= "10000101"; x_in <= "00001010"; z_correct<="1111101100110010";
        when 1419 => y_in <= "10000101"; x_in <= "00001011"; z_correct<="1111101010110111";
        when 1420 => y_in <= "10000101"; x_in <= "00001100"; z_correct<="1111101000111100";
        when 1421 => y_in <= "10000101"; x_in <= "00001101"; z_correct<="1111100111000001";
        when 1422 => y_in <= "10000101"; x_in <= "00001110"; z_correct<="1111100101000110";
        when 1423 => y_in <= "10000101"; x_in <= "00001111"; z_correct<="1111100011001011";
        when 1424 => y_in <= "10000101"; x_in <= "00010000"; z_correct<="1111100001010000";
        when 1425 => y_in <= "10000101"; x_in <= "00010001"; z_correct<="1111011111010101";
        when 1426 => y_in <= "10000101"; x_in <= "00010010"; z_correct<="1111011101011010";
        when 1427 => y_in <= "10000101"; x_in <= "00010011"; z_correct<="1111011011011111";
        when 1428 => y_in <= "10000101"; x_in <= "00010100"; z_correct<="1111011001100100";
        when 1429 => y_in <= "10000101"; x_in <= "00010101"; z_correct<="1111010111101001";
        when 1430 => y_in <= "10000101"; x_in <= "00010110"; z_correct<="1111010101101110";
        when 1431 => y_in <= "10000101"; x_in <= "00010111"; z_correct<="1111010011110011";
        when 1432 => y_in <= "10000101"; x_in <= "00011000"; z_correct<="1111010001111000";
        when 1433 => y_in <= "10000101"; x_in <= "00011001"; z_correct<="1111001111111101";
        when 1434 => y_in <= "10000101"; x_in <= "00011010"; z_correct<="1111001110000010";
        when 1435 => y_in <= "10000101"; x_in <= "00011011"; z_correct<="1111001100000111";
        when 1436 => y_in <= "10000101"; x_in <= "00011100"; z_correct<="1111001010001100";
        when 1437 => y_in <= "10000101"; x_in <= "00011101"; z_correct<="1111001000010001";
        when 1438 => y_in <= "10000101"; x_in <= "00011110"; z_correct<="1111000110010110";
        when 1439 => y_in <= "10000101"; x_in <= "00011111"; z_correct<="1111000100011011";
        when 1440 => y_in <= "10000101"; x_in <= "00100000"; z_correct<="1111000010100000";
        when 1441 => y_in <= "10000101"; x_in <= "00100001"; z_correct<="1111000000100101";
        when 1442 => y_in <= "10000101"; x_in <= "00100010"; z_correct<="1110111110101010";
        when 1443 => y_in <= "10000101"; x_in <= "00100011"; z_correct<="1110111100101111";
        when 1444 => y_in <= "10000101"; x_in <= "00100100"; z_correct<="1110111010110100";
        when 1445 => y_in <= "10000101"; x_in <= "00100101"; z_correct<="1110111000111001";
        when 1446 => y_in <= "10000101"; x_in <= "00100110"; z_correct<="1110110110111110";
        when 1447 => y_in <= "10000101"; x_in <= "00100111"; z_correct<="1110110101000011";
        when 1448 => y_in <= "10000101"; x_in <= "00101000"; z_correct<="1110110011001000";
        when 1449 => y_in <= "10000101"; x_in <= "00101001"; z_correct<="1110110001001101";
        when 1450 => y_in <= "10000101"; x_in <= "00101010"; z_correct<="1110101111010010";
        when 1451 => y_in <= "10000101"; x_in <= "00101011"; z_correct<="1110101101010111";
        when 1452 => y_in <= "10000101"; x_in <= "00101100"; z_correct<="1110101011011100";
        when 1453 => y_in <= "10000101"; x_in <= "00101101"; z_correct<="1110101001100001";
        when 1454 => y_in <= "10000101"; x_in <= "00101110"; z_correct<="1110100111100110";
        when 1455 => y_in <= "10000101"; x_in <= "00101111"; z_correct<="1110100101101011";
        when 1456 => y_in <= "10000101"; x_in <= "00110000"; z_correct<="1110100011110000";
        when 1457 => y_in <= "10000101"; x_in <= "00110001"; z_correct<="1110100001110101";
        when 1458 => y_in <= "10000101"; x_in <= "00110010"; z_correct<="1110011111111010";
        when 1459 => y_in <= "10000101"; x_in <= "00110011"; z_correct<="1110011101111111";
        when 1460 => y_in <= "10000101"; x_in <= "00110100"; z_correct<="1110011100000100";
        when 1461 => y_in <= "10000101"; x_in <= "00110101"; z_correct<="1110011010001001";
        when 1462 => y_in <= "10000101"; x_in <= "00110110"; z_correct<="1110011000001110";
        when 1463 => y_in <= "10000101"; x_in <= "00110111"; z_correct<="1110010110010011";
        when 1464 => y_in <= "10000101"; x_in <= "00111000"; z_correct<="1110010100011000";
        when 1465 => y_in <= "10000101"; x_in <= "00111001"; z_correct<="1110010010011101";
        when 1466 => y_in <= "10000101"; x_in <= "00111010"; z_correct<="1110010000100010";
        when 1467 => y_in <= "10000101"; x_in <= "00111011"; z_correct<="1110001110100111";
        when 1468 => y_in <= "10000101"; x_in <= "00111100"; z_correct<="1110001100101100";
        when 1469 => y_in <= "10000101"; x_in <= "00111101"; z_correct<="1110001010110001";
        when 1470 => y_in <= "10000101"; x_in <= "00111110"; z_correct<="1110001000110110";
        when 1471 => y_in <= "10000101"; x_in <= "00111111"; z_correct<="1110000110111011";
        when 1472 => y_in <= "10000101"; x_in <= "01000000"; z_correct<="1110000101000000";
        when 1473 => y_in <= "10000101"; x_in <= "01000001"; z_correct<="1110000011000101";
        when 1474 => y_in <= "10000101"; x_in <= "01000010"; z_correct<="1110000001001010";
        when 1475 => y_in <= "10000101"; x_in <= "01000011"; z_correct<="1101111111001111";
        when 1476 => y_in <= "10000101"; x_in <= "01000100"; z_correct<="1101111101010100";
        when 1477 => y_in <= "10000101"; x_in <= "01000101"; z_correct<="1101111011011001";
        when 1478 => y_in <= "10000101"; x_in <= "01000110"; z_correct<="1101111001011110";
        when 1479 => y_in <= "10000101"; x_in <= "01000111"; z_correct<="1101110111100011";
        when 1480 => y_in <= "10000101"; x_in <= "01001000"; z_correct<="1101110101101000";
        when 1481 => y_in <= "10000101"; x_in <= "01001001"; z_correct<="1101110011101101";
        when 1482 => y_in <= "10000101"; x_in <= "01001010"; z_correct<="1101110001110010";
        when 1483 => y_in <= "10000101"; x_in <= "01001011"; z_correct<="1101101111110111";
        when 1484 => y_in <= "10000101"; x_in <= "01001100"; z_correct<="1101101101111100";
        when 1485 => y_in <= "10000101"; x_in <= "01001101"; z_correct<="1101101100000001";
        when 1486 => y_in <= "10000101"; x_in <= "01001110"; z_correct<="1101101010000110";
        when 1487 => y_in <= "10000101"; x_in <= "01001111"; z_correct<="1101101000001011";
        when 1488 => y_in <= "10000101"; x_in <= "01010000"; z_correct<="1101100110010000";
        when 1489 => y_in <= "10000101"; x_in <= "01010001"; z_correct<="1101100100010101";
        when 1490 => y_in <= "10000101"; x_in <= "01010010"; z_correct<="1101100010011010";
        when 1491 => y_in <= "10000101"; x_in <= "01010011"; z_correct<="1101100000011111";
        when 1492 => y_in <= "10000101"; x_in <= "01010100"; z_correct<="1101011110100100";
        when 1493 => y_in <= "10000101"; x_in <= "01010101"; z_correct<="1101011100101001";
        when 1494 => y_in <= "10000101"; x_in <= "01010110"; z_correct<="1101011010101110";
        when 1495 => y_in <= "10000101"; x_in <= "01010111"; z_correct<="1101011000110011";
        when 1496 => y_in <= "10000101"; x_in <= "01011000"; z_correct<="1101010110111000";
        when 1497 => y_in <= "10000101"; x_in <= "01011001"; z_correct<="1101010100111101";
        when 1498 => y_in <= "10000101"; x_in <= "01011010"; z_correct<="1101010011000010";
        when 1499 => y_in <= "10000101"; x_in <= "01011011"; z_correct<="1101010001000111";
        when 1500 => y_in <= "10000101"; x_in <= "01011100"; z_correct<="1101001111001100";
        when 1501 => y_in <= "10000101"; x_in <= "01011101"; z_correct<="1101001101010001";
        when 1502 => y_in <= "10000101"; x_in <= "01011110"; z_correct<="1101001011010110";
        when 1503 => y_in <= "10000101"; x_in <= "01011111"; z_correct<="1101001001011011";
        when 1504 => y_in <= "10000101"; x_in <= "01100000"; z_correct<="1101000111100000";
        when 1505 => y_in <= "10000101"; x_in <= "01100001"; z_correct<="1101000101100101";
        when 1506 => y_in <= "10000101"; x_in <= "01100010"; z_correct<="1101000011101010";
        when 1507 => y_in <= "10000101"; x_in <= "01100011"; z_correct<="1101000001101111";
        when 1508 => y_in <= "10000101"; x_in <= "01100100"; z_correct<="1100111111110100";
        when 1509 => y_in <= "10000101"; x_in <= "01100101"; z_correct<="1100111101111001";
        when 1510 => y_in <= "10000101"; x_in <= "01100110"; z_correct<="1100111011111110";
        when 1511 => y_in <= "10000101"; x_in <= "01100111"; z_correct<="1100111010000011";
        when 1512 => y_in <= "10000101"; x_in <= "01101000"; z_correct<="1100111000001000";
        when 1513 => y_in <= "10000101"; x_in <= "01101001"; z_correct<="1100110110001101";
        when 1514 => y_in <= "10000101"; x_in <= "01101010"; z_correct<="1100110100010010";
        when 1515 => y_in <= "10000101"; x_in <= "01101011"; z_correct<="1100110010010111";
        when 1516 => y_in <= "10000101"; x_in <= "01101100"; z_correct<="1100110000011100";
        when 1517 => y_in <= "10000101"; x_in <= "01101101"; z_correct<="1100101110100001";
        when 1518 => y_in <= "10000101"; x_in <= "01101110"; z_correct<="1100101100100110";
        when 1519 => y_in <= "10000101"; x_in <= "01101111"; z_correct<="1100101010101011";
        when 1520 => y_in <= "10000101"; x_in <= "01110000"; z_correct<="1100101000110000";
        when 1521 => y_in <= "10000101"; x_in <= "01110001"; z_correct<="1100100110110101";
        when 1522 => y_in <= "10000101"; x_in <= "01110010"; z_correct<="1100100100111010";
        when 1523 => y_in <= "10000101"; x_in <= "01110011"; z_correct<="1100100010111111";
        when 1524 => y_in <= "10000101"; x_in <= "01110100"; z_correct<="1100100001000100";
        when 1525 => y_in <= "10000101"; x_in <= "01110101"; z_correct<="1100011111001001";
        when 1526 => y_in <= "10000101"; x_in <= "01110110"; z_correct<="1100011101001110";
        when 1527 => y_in <= "10000101"; x_in <= "01110111"; z_correct<="1100011011010011";
        when 1528 => y_in <= "10000101"; x_in <= "01111000"; z_correct<="1100011001011000";
        when 1529 => y_in <= "10000101"; x_in <= "01111001"; z_correct<="1100010111011101";
        when 1530 => y_in <= "10000101"; x_in <= "01111010"; z_correct<="1100010101100010";
        when 1531 => y_in <= "10000101"; x_in <= "01111011"; z_correct<="1100010011100111";
        when 1532 => y_in <= "10000101"; x_in <= "01111100"; z_correct<="1100010001101100";
        when 1533 => y_in <= "10000101"; x_in <= "01111101"; z_correct<="1100001111110001";
        when 1534 => y_in <= "10000101"; x_in <= "01111110"; z_correct<="1100001101110110";
        when 1535 => y_in <= "10000101"; x_in <= "01111111"; z_correct<="1100001011111011";
        when 1536 => y_in <= "10000110"; x_in <= "10000000"; z_correct<="0011110100000000";
        when 1537 => y_in <= "10000110"; x_in <= "10000001"; z_correct<="0011110010000110";
        when 1538 => y_in <= "10000110"; x_in <= "10000010"; z_correct<="0011110000001100";
        when 1539 => y_in <= "10000110"; x_in <= "10000011"; z_correct<="0011101110010010";
        when 1540 => y_in <= "10000110"; x_in <= "10000100"; z_correct<="0011101100011000";
        when 1541 => y_in <= "10000110"; x_in <= "10000101"; z_correct<="0011101010011110";
        when 1542 => y_in <= "10000110"; x_in <= "10000110"; z_correct<="0011101000100100";
        when 1543 => y_in <= "10000110"; x_in <= "10000111"; z_correct<="0011100110101010";
        when 1544 => y_in <= "10000110"; x_in <= "10001000"; z_correct<="0011100100110000";
        when 1545 => y_in <= "10000110"; x_in <= "10001001"; z_correct<="0011100010110110";
        when 1546 => y_in <= "10000110"; x_in <= "10001010"; z_correct<="0011100000111100";
        when 1547 => y_in <= "10000110"; x_in <= "10001011"; z_correct<="0011011111000010";
        when 1548 => y_in <= "10000110"; x_in <= "10001100"; z_correct<="0011011101001000";
        when 1549 => y_in <= "10000110"; x_in <= "10001101"; z_correct<="0011011011001110";
        when 1550 => y_in <= "10000110"; x_in <= "10001110"; z_correct<="0011011001010100";
        when 1551 => y_in <= "10000110"; x_in <= "10001111"; z_correct<="0011010111011010";
        when 1552 => y_in <= "10000110"; x_in <= "10010000"; z_correct<="0011010101100000";
        when 1553 => y_in <= "10000110"; x_in <= "10010001"; z_correct<="0011010011100110";
        when 1554 => y_in <= "10000110"; x_in <= "10010010"; z_correct<="0011010001101100";
        when 1555 => y_in <= "10000110"; x_in <= "10010011"; z_correct<="0011001111110010";
        when 1556 => y_in <= "10000110"; x_in <= "10010100"; z_correct<="0011001101111000";
        when 1557 => y_in <= "10000110"; x_in <= "10010101"; z_correct<="0011001011111110";
        when 1558 => y_in <= "10000110"; x_in <= "10010110"; z_correct<="0011001010000100";
        when 1559 => y_in <= "10000110"; x_in <= "10010111"; z_correct<="0011001000001010";
        when 1560 => y_in <= "10000110"; x_in <= "10011000"; z_correct<="0011000110010000";
        when 1561 => y_in <= "10000110"; x_in <= "10011001"; z_correct<="0011000100010110";
        when 1562 => y_in <= "10000110"; x_in <= "10011010"; z_correct<="0011000010011100";
        when 1563 => y_in <= "10000110"; x_in <= "10011011"; z_correct<="0011000000100010";
        when 1564 => y_in <= "10000110"; x_in <= "10011100"; z_correct<="0010111110101000";
        when 1565 => y_in <= "10000110"; x_in <= "10011101"; z_correct<="0010111100101110";
        when 1566 => y_in <= "10000110"; x_in <= "10011110"; z_correct<="0010111010110100";
        when 1567 => y_in <= "10000110"; x_in <= "10011111"; z_correct<="0010111000111010";
        when 1568 => y_in <= "10000110"; x_in <= "10100000"; z_correct<="0010110111000000";
        when 1569 => y_in <= "10000110"; x_in <= "10100001"; z_correct<="0010110101000110";
        when 1570 => y_in <= "10000110"; x_in <= "10100010"; z_correct<="0010110011001100";
        when 1571 => y_in <= "10000110"; x_in <= "10100011"; z_correct<="0010110001010010";
        when 1572 => y_in <= "10000110"; x_in <= "10100100"; z_correct<="0010101111011000";
        when 1573 => y_in <= "10000110"; x_in <= "10100101"; z_correct<="0010101101011110";
        when 1574 => y_in <= "10000110"; x_in <= "10100110"; z_correct<="0010101011100100";
        when 1575 => y_in <= "10000110"; x_in <= "10100111"; z_correct<="0010101001101010";
        when 1576 => y_in <= "10000110"; x_in <= "10101000"; z_correct<="0010100111110000";
        when 1577 => y_in <= "10000110"; x_in <= "10101001"; z_correct<="0010100101110110";
        when 1578 => y_in <= "10000110"; x_in <= "10101010"; z_correct<="0010100011111100";
        when 1579 => y_in <= "10000110"; x_in <= "10101011"; z_correct<="0010100010000010";
        when 1580 => y_in <= "10000110"; x_in <= "10101100"; z_correct<="0010100000001000";
        when 1581 => y_in <= "10000110"; x_in <= "10101101"; z_correct<="0010011110001110";
        when 1582 => y_in <= "10000110"; x_in <= "10101110"; z_correct<="0010011100010100";
        when 1583 => y_in <= "10000110"; x_in <= "10101111"; z_correct<="0010011010011010";
        when 1584 => y_in <= "10000110"; x_in <= "10110000"; z_correct<="0010011000100000";
        when 1585 => y_in <= "10000110"; x_in <= "10110001"; z_correct<="0010010110100110";
        when 1586 => y_in <= "10000110"; x_in <= "10110010"; z_correct<="0010010100101100";
        when 1587 => y_in <= "10000110"; x_in <= "10110011"; z_correct<="0010010010110010";
        when 1588 => y_in <= "10000110"; x_in <= "10110100"; z_correct<="0010010000111000";
        when 1589 => y_in <= "10000110"; x_in <= "10110101"; z_correct<="0010001110111110";
        when 1590 => y_in <= "10000110"; x_in <= "10110110"; z_correct<="0010001101000100";
        when 1591 => y_in <= "10000110"; x_in <= "10110111"; z_correct<="0010001011001010";
        when 1592 => y_in <= "10000110"; x_in <= "10111000"; z_correct<="0010001001010000";
        when 1593 => y_in <= "10000110"; x_in <= "10111001"; z_correct<="0010000111010110";
        when 1594 => y_in <= "10000110"; x_in <= "10111010"; z_correct<="0010000101011100";
        when 1595 => y_in <= "10000110"; x_in <= "10111011"; z_correct<="0010000011100010";
        when 1596 => y_in <= "10000110"; x_in <= "10111100"; z_correct<="0010000001101000";
        when 1597 => y_in <= "10000110"; x_in <= "10111101"; z_correct<="0001111111101110";
        when 1598 => y_in <= "10000110"; x_in <= "10111110"; z_correct<="0001111101110100";
        when 1599 => y_in <= "10000110"; x_in <= "10111111"; z_correct<="0001111011111010";
        when 1600 => y_in <= "10000110"; x_in <= "11000000"; z_correct<="0001111010000000";
        when 1601 => y_in <= "10000110"; x_in <= "11000001"; z_correct<="0001111000000110";
        when 1602 => y_in <= "10000110"; x_in <= "11000010"; z_correct<="0001110110001100";
        when 1603 => y_in <= "10000110"; x_in <= "11000011"; z_correct<="0001110100010010";
        when 1604 => y_in <= "10000110"; x_in <= "11000100"; z_correct<="0001110010011000";
        when 1605 => y_in <= "10000110"; x_in <= "11000101"; z_correct<="0001110000011110";
        when 1606 => y_in <= "10000110"; x_in <= "11000110"; z_correct<="0001101110100100";
        when 1607 => y_in <= "10000110"; x_in <= "11000111"; z_correct<="0001101100101010";
        when 1608 => y_in <= "10000110"; x_in <= "11001000"; z_correct<="0001101010110000";
        when 1609 => y_in <= "10000110"; x_in <= "11001001"; z_correct<="0001101000110110";
        when 1610 => y_in <= "10000110"; x_in <= "11001010"; z_correct<="0001100110111100";
        when 1611 => y_in <= "10000110"; x_in <= "11001011"; z_correct<="0001100101000010";
        when 1612 => y_in <= "10000110"; x_in <= "11001100"; z_correct<="0001100011001000";
        when 1613 => y_in <= "10000110"; x_in <= "11001101"; z_correct<="0001100001001110";
        when 1614 => y_in <= "10000110"; x_in <= "11001110"; z_correct<="0001011111010100";
        when 1615 => y_in <= "10000110"; x_in <= "11001111"; z_correct<="0001011101011010";
        when 1616 => y_in <= "10000110"; x_in <= "11010000"; z_correct<="0001011011100000";
        when 1617 => y_in <= "10000110"; x_in <= "11010001"; z_correct<="0001011001100110";
        when 1618 => y_in <= "10000110"; x_in <= "11010010"; z_correct<="0001010111101100";
        when 1619 => y_in <= "10000110"; x_in <= "11010011"; z_correct<="0001010101110010";
        when 1620 => y_in <= "10000110"; x_in <= "11010100"; z_correct<="0001010011111000";
        when 1621 => y_in <= "10000110"; x_in <= "11010101"; z_correct<="0001010001111110";
        when 1622 => y_in <= "10000110"; x_in <= "11010110"; z_correct<="0001010000000100";
        when 1623 => y_in <= "10000110"; x_in <= "11010111"; z_correct<="0001001110001010";
        when 1624 => y_in <= "10000110"; x_in <= "11011000"; z_correct<="0001001100010000";
        when 1625 => y_in <= "10000110"; x_in <= "11011001"; z_correct<="0001001010010110";
        when 1626 => y_in <= "10000110"; x_in <= "11011010"; z_correct<="0001001000011100";
        when 1627 => y_in <= "10000110"; x_in <= "11011011"; z_correct<="0001000110100010";
        when 1628 => y_in <= "10000110"; x_in <= "11011100"; z_correct<="0001000100101000";
        when 1629 => y_in <= "10000110"; x_in <= "11011101"; z_correct<="0001000010101110";
        when 1630 => y_in <= "10000110"; x_in <= "11011110"; z_correct<="0001000000110100";
        when 1631 => y_in <= "10000110"; x_in <= "11011111"; z_correct<="0000111110111010";
        when 1632 => y_in <= "10000110"; x_in <= "11100000"; z_correct<="0000111101000000";
        when 1633 => y_in <= "10000110"; x_in <= "11100001"; z_correct<="0000111011000110";
        when 1634 => y_in <= "10000110"; x_in <= "11100010"; z_correct<="0000111001001100";
        when 1635 => y_in <= "10000110"; x_in <= "11100011"; z_correct<="0000110111010010";
        when 1636 => y_in <= "10000110"; x_in <= "11100100"; z_correct<="0000110101011000";
        when 1637 => y_in <= "10000110"; x_in <= "11100101"; z_correct<="0000110011011110";
        when 1638 => y_in <= "10000110"; x_in <= "11100110"; z_correct<="0000110001100100";
        when 1639 => y_in <= "10000110"; x_in <= "11100111"; z_correct<="0000101111101010";
        when 1640 => y_in <= "10000110"; x_in <= "11101000"; z_correct<="0000101101110000";
        when 1641 => y_in <= "10000110"; x_in <= "11101001"; z_correct<="0000101011110110";
        when 1642 => y_in <= "10000110"; x_in <= "11101010"; z_correct<="0000101001111100";
        when 1643 => y_in <= "10000110"; x_in <= "11101011"; z_correct<="0000101000000010";
        when 1644 => y_in <= "10000110"; x_in <= "11101100"; z_correct<="0000100110001000";
        when 1645 => y_in <= "10000110"; x_in <= "11101101"; z_correct<="0000100100001110";
        when 1646 => y_in <= "10000110"; x_in <= "11101110"; z_correct<="0000100010010100";
        when 1647 => y_in <= "10000110"; x_in <= "11101111"; z_correct<="0000100000011010";
        when 1648 => y_in <= "10000110"; x_in <= "11110000"; z_correct<="0000011110100000";
        when 1649 => y_in <= "10000110"; x_in <= "11110001"; z_correct<="0000011100100110";
        when 1650 => y_in <= "10000110"; x_in <= "11110010"; z_correct<="0000011010101100";
        when 1651 => y_in <= "10000110"; x_in <= "11110011"; z_correct<="0000011000110010";
        when 1652 => y_in <= "10000110"; x_in <= "11110100"; z_correct<="0000010110111000";
        when 1653 => y_in <= "10000110"; x_in <= "11110101"; z_correct<="0000010100111110";
        when 1654 => y_in <= "10000110"; x_in <= "11110110"; z_correct<="0000010011000100";
        when 1655 => y_in <= "10000110"; x_in <= "11110111"; z_correct<="0000010001001010";
        when 1656 => y_in <= "10000110"; x_in <= "11111000"; z_correct<="0000001111010000";
        when 1657 => y_in <= "10000110"; x_in <= "11111001"; z_correct<="0000001101010110";
        when 1658 => y_in <= "10000110"; x_in <= "11111010"; z_correct<="0000001011011100";
        when 1659 => y_in <= "10000110"; x_in <= "11111011"; z_correct<="0000001001100010";
        when 1660 => y_in <= "10000110"; x_in <= "11111100"; z_correct<="0000000111101000";
        when 1661 => y_in <= "10000110"; x_in <= "11111101"; z_correct<="0000000101101110";
        when 1662 => y_in <= "10000110"; x_in <= "11111110"; z_correct<="0000000011110100";
        when 1663 => y_in <= "10000110"; x_in <= "11111111"; z_correct<="0000000001111010";
        when 1664 => y_in <= "10000110"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 1665 => y_in <= "10000110"; x_in <= "00000001"; z_correct<="1111111110000110";
        when 1666 => y_in <= "10000110"; x_in <= "00000010"; z_correct<="1111111100001100";
        when 1667 => y_in <= "10000110"; x_in <= "00000011"; z_correct<="1111111010010010";
        when 1668 => y_in <= "10000110"; x_in <= "00000100"; z_correct<="1111111000011000";
        when 1669 => y_in <= "10000110"; x_in <= "00000101"; z_correct<="1111110110011110";
        when 1670 => y_in <= "10000110"; x_in <= "00000110"; z_correct<="1111110100100100";
        when 1671 => y_in <= "10000110"; x_in <= "00000111"; z_correct<="1111110010101010";
        when 1672 => y_in <= "10000110"; x_in <= "00001000"; z_correct<="1111110000110000";
        when 1673 => y_in <= "10000110"; x_in <= "00001001"; z_correct<="1111101110110110";
        when 1674 => y_in <= "10000110"; x_in <= "00001010"; z_correct<="1111101100111100";
        when 1675 => y_in <= "10000110"; x_in <= "00001011"; z_correct<="1111101011000010";
        when 1676 => y_in <= "10000110"; x_in <= "00001100"; z_correct<="1111101001001000";
        when 1677 => y_in <= "10000110"; x_in <= "00001101"; z_correct<="1111100111001110";
        when 1678 => y_in <= "10000110"; x_in <= "00001110"; z_correct<="1111100101010100";
        when 1679 => y_in <= "10000110"; x_in <= "00001111"; z_correct<="1111100011011010";
        when 1680 => y_in <= "10000110"; x_in <= "00010000"; z_correct<="1111100001100000";
        when 1681 => y_in <= "10000110"; x_in <= "00010001"; z_correct<="1111011111100110";
        when 1682 => y_in <= "10000110"; x_in <= "00010010"; z_correct<="1111011101101100";
        when 1683 => y_in <= "10000110"; x_in <= "00010011"; z_correct<="1111011011110010";
        when 1684 => y_in <= "10000110"; x_in <= "00010100"; z_correct<="1111011001111000";
        when 1685 => y_in <= "10000110"; x_in <= "00010101"; z_correct<="1111010111111110";
        when 1686 => y_in <= "10000110"; x_in <= "00010110"; z_correct<="1111010110000100";
        when 1687 => y_in <= "10000110"; x_in <= "00010111"; z_correct<="1111010100001010";
        when 1688 => y_in <= "10000110"; x_in <= "00011000"; z_correct<="1111010010010000";
        when 1689 => y_in <= "10000110"; x_in <= "00011001"; z_correct<="1111010000010110";
        when 1690 => y_in <= "10000110"; x_in <= "00011010"; z_correct<="1111001110011100";
        when 1691 => y_in <= "10000110"; x_in <= "00011011"; z_correct<="1111001100100010";
        when 1692 => y_in <= "10000110"; x_in <= "00011100"; z_correct<="1111001010101000";
        when 1693 => y_in <= "10000110"; x_in <= "00011101"; z_correct<="1111001000101110";
        when 1694 => y_in <= "10000110"; x_in <= "00011110"; z_correct<="1111000110110100";
        when 1695 => y_in <= "10000110"; x_in <= "00011111"; z_correct<="1111000100111010";
        when 1696 => y_in <= "10000110"; x_in <= "00100000"; z_correct<="1111000011000000";
        when 1697 => y_in <= "10000110"; x_in <= "00100001"; z_correct<="1111000001000110";
        when 1698 => y_in <= "10000110"; x_in <= "00100010"; z_correct<="1110111111001100";
        when 1699 => y_in <= "10000110"; x_in <= "00100011"; z_correct<="1110111101010010";
        when 1700 => y_in <= "10000110"; x_in <= "00100100"; z_correct<="1110111011011000";
        when 1701 => y_in <= "10000110"; x_in <= "00100101"; z_correct<="1110111001011110";
        when 1702 => y_in <= "10000110"; x_in <= "00100110"; z_correct<="1110110111100100";
        when 1703 => y_in <= "10000110"; x_in <= "00100111"; z_correct<="1110110101101010";
        when 1704 => y_in <= "10000110"; x_in <= "00101000"; z_correct<="1110110011110000";
        when 1705 => y_in <= "10000110"; x_in <= "00101001"; z_correct<="1110110001110110";
        when 1706 => y_in <= "10000110"; x_in <= "00101010"; z_correct<="1110101111111100";
        when 1707 => y_in <= "10000110"; x_in <= "00101011"; z_correct<="1110101110000010";
        when 1708 => y_in <= "10000110"; x_in <= "00101100"; z_correct<="1110101100001000";
        when 1709 => y_in <= "10000110"; x_in <= "00101101"; z_correct<="1110101010001110";
        when 1710 => y_in <= "10000110"; x_in <= "00101110"; z_correct<="1110101000010100";
        when 1711 => y_in <= "10000110"; x_in <= "00101111"; z_correct<="1110100110011010";
        when 1712 => y_in <= "10000110"; x_in <= "00110000"; z_correct<="1110100100100000";
        when 1713 => y_in <= "10000110"; x_in <= "00110001"; z_correct<="1110100010100110";
        when 1714 => y_in <= "10000110"; x_in <= "00110010"; z_correct<="1110100000101100";
        when 1715 => y_in <= "10000110"; x_in <= "00110011"; z_correct<="1110011110110010";
        when 1716 => y_in <= "10000110"; x_in <= "00110100"; z_correct<="1110011100111000";
        when 1717 => y_in <= "10000110"; x_in <= "00110101"; z_correct<="1110011010111110";
        when 1718 => y_in <= "10000110"; x_in <= "00110110"; z_correct<="1110011001000100";
        when 1719 => y_in <= "10000110"; x_in <= "00110111"; z_correct<="1110010111001010";
        when 1720 => y_in <= "10000110"; x_in <= "00111000"; z_correct<="1110010101010000";
        when 1721 => y_in <= "10000110"; x_in <= "00111001"; z_correct<="1110010011010110";
        when 1722 => y_in <= "10000110"; x_in <= "00111010"; z_correct<="1110010001011100";
        when 1723 => y_in <= "10000110"; x_in <= "00111011"; z_correct<="1110001111100010";
        when 1724 => y_in <= "10000110"; x_in <= "00111100"; z_correct<="1110001101101000";
        when 1725 => y_in <= "10000110"; x_in <= "00111101"; z_correct<="1110001011101110";
        when 1726 => y_in <= "10000110"; x_in <= "00111110"; z_correct<="1110001001110100";
        when 1727 => y_in <= "10000110"; x_in <= "00111111"; z_correct<="1110000111111010";
        when 1728 => y_in <= "10000110"; x_in <= "01000000"; z_correct<="1110000110000000";
        when 1729 => y_in <= "10000110"; x_in <= "01000001"; z_correct<="1110000100000110";
        when 1730 => y_in <= "10000110"; x_in <= "01000010"; z_correct<="1110000010001100";
        when 1731 => y_in <= "10000110"; x_in <= "01000011"; z_correct<="1110000000010010";
        when 1732 => y_in <= "10000110"; x_in <= "01000100"; z_correct<="1101111110011000";
        when 1733 => y_in <= "10000110"; x_in <= "01000101"; z_correct<="1101111100011110";
        when 1734 => y_in <= "10000110"; x_in <= "01000110"; z_correct<="1101111010100100";
        when 1735 => y_in <= "10000110"; x_in <= "01000111"; z_correct<="1101111000101010";
        when 1736 => y_in <= "10000110"; x_in <= "01001000"; z_correct<="1101110110110000";
        when 1737 => y_in <= "10000110"; x_in <= "01001001"; z_correct<="1101110100110110";
        when 1738 => y_in <= "10000110"; x_in <= "01001010"; z_correct<="1101110010111100";
        when 1739 => y_in <= "10000110"; x_in <= "01001011"; z_correct<="1101110001000010";
        when 1740 => y_in <= "10000110"; x_in <= "01001100"; z_correct<="1101101111001000";
        when 1741 => y_in <= "10000110"; x_in <= "01001101"; z_correct<="1101101101001110";
        when 1742 => y_in <= "10000110"; x_in <= "01001110"; z_correct<="1101101011010100";
        when 1743 => y_in <= "10000110"; x_in <= "01001111"; z_correct<="1101101001011010";
        when 1744 => y_in <= "10000110"; x_in <= "01010000"; z_correct<="1101100111100000";
        when 1745 => y_in <= "10000110"; x_in <= "01010001"; z_correct<="1101100101100110";
        when 1746 => y_in <= "10000110"; x_in <= "01010010"; z_correct<="1101100011101100";
        when 1747 => y_in <= "10000110"; x_in <= "01010011"; z_correct<="1101100001110010";
        when 1748 => y_in <= "10000110"; x_in <= "01010100"; z_correct<="1101011111111000";
        when 1749 => y_in <= "10000110"; x_in <= "01010101"; z_correct<="1101011101111110";
        when 1750 => y_in <= "10000110"; x_in <= "01010110"; z_correct<="1101011100000100";
        when 1751 => y_in <= "10000110"; x_in <= "01010111"; z_correct<="1101011010001010";
        when 1752 => y_in <= "10000110"; x_in <= "01011000"; z_correct<="1101011000010000";
        when 1753 => y_in <= "10000110"; x_in <= "01011001"; z_correct<="1101010110010110";
        when 1754 => y_in <= "10000110"; x_in <= "01011010"; z_correct<="1101010100011100";
        when 1755 => y_in <= "10000110"; x_in <= "01011011"; z_correct<="1101010010100010";
        when 1756 => y_in <= "10000110"; x_in <= "01011100"; z_correct<="1101010000101000";
        when 1757 => y_in <= "10000110"; x_in <= "01011101"; z_correct<="1101001110101110";
        when 1758 => y_in <= "10000110"; x_in <= "01011110"; z_correct<="1101001100110100";
        when 1759 => y_in <= "10000110"; x_in <= "01011111"; z_correct<="1101001010111010";
        when 1760 => y_in <= "10000110"; x_in <= "01100000"; z_correct<="1101001001000000";
        when 1761 => y_in <= "10000110"; x_in <= "01100001"; z_correct<="1101000111000110";
        when 1762 => y_in <= "10000110"; x_in <= "01100010"; z_correct<="1101000101001100";
        when 1763 => y_in <= "10000110"; x_in <= "01100011"; z_correct<="1101000011010010";
        when 1764 => y_in <= "10000110"; x_in <= "01100100"; z_correct<="1101000001011000";
        when 1765 => y_in <= "10000110"; x_in <= "01100101"; z_correct<="1100111111011110";
        when 1766 => y_in <= "10000110"; x_in <= "01100110"; z_correct<="1100111101100100";
        when 1767 => y_in <= "10000110"; x_in <= "01100111"; z_correct<="1100111011101010";
        when 1768 => y_in <= "10000110"; x_in <= "01101000"; z_correct<="1100111001110000";
        when 1769 => y_in <= "10000110"; x_in <= "01101001"; z_correct<="1100110111110110";
        when 1770 => y_in <= "10000110"; x_in <= "01101010"; z_correct<="1100110101111100";
        when 1771 => y_in <= "10000110"; x_in <= "01101011"; z_correct<="1100110100000010";
        when 1772 => y_in <= "10000110"; x_in <= "01101100"; z_correct<="1100110010001000";
        when 1773 => y_in <= "10000110"; x_in <= "01101101"; z_correct<="1100110000001110";
        when 1774 => y_in <= "10000110"; x_in <= "01101110"; z_correct<="1100101110010100";
        when 1775 => y_in <= "10000110"; x_in <= "01101111"; z_correct<="1100101100011010";
        when 1776 => y_in <= "10000110"; x_in <= "01110000"; z_correct<="1100101010100000";
        when 1777 => y_in <= "10000110"; x_in <= "01110001"; z_correct<="1100101000100110";
        when 1778 => y_in <= "10000110"; x_in <= "01110010"; z_correct<="1100100110101100";
        when 1779 => y_in <= "10000110"; x_in <= "01110011"; z_correct<="1100100100110010";
        when 1780 => y_in <= "10000110"; x_in <= "01110100"; z_correct<="1100100010111000";
        when 1781 => y_in <= "10000110"; x_in <= "01110101"; z_correct<="1100100000111110";
        when 1782 => y_in <= "10000110"; x_in <= "01110110"; z_correct<="1100011111000100";
        when 1783 => y_in <= "10000110"; x_in <= "01110111"; z_correct<="1100011101001010";
        when 1784 => y_in <= "10000110"; x_in <= "01111000"; z_correct<="1100011011010000";
        when 1785 => y_in <= "10000110"; x_in <= "01111001"; z_correct<="1100011001010110";
        when 1786 => y_in <= "10000110"; x_in <= "01111010"; z_correct<="1100010111011100";
        when 1787 => y_in <= "10000110"; x_in <= "01111011"; z_correct<="1100010101100010";
        when 1788 => y_in <= "10000110"; x_in <= "01111100"; z_correct<="1100010011101000";
        when 1789 => y_in <= "10000110"; x_in <= "01111101"; z_correct<="1100010001101110";
        when 1790 => y_in <= "10000110"; x_in <= "01111110"; z_correct<="1100001111110100";
        when 1791 => y_in <= "10000110"; x_in <= "01111111"; z_correct<="1100001101111010";
        when 1792 => y_in <= "10000111"; x_in <= "10000000"; z_correct<="0011110010000000";
        when 1793 => y_in <= "10000111"; x_in <= "10000001"; z_correct<="0011110000000111";
        when 1794 => y_in <= "10000111"; x_in <= "10000010"; z_correct<="0011101110001110";
        when 1795 => y_in <= "10000111"; x_in <= "10000011"; z_correct<="0011101100010101";
        when 1796 => y_in <= "10000111"; x_in <= "10000100"; z_correct<="0011101010011100";
        when 1797 => y_in <= "10000111"; x_in <= "10000101"; z_correct<="0011101000100011";
        when 1798 => y_in <= "10000111"; x_in <= "10000110"; z_correct<="0011100110101010";
        when 1799 => y_in <= "10000111"; x_in <= "10000111"; z_correct<="0011100100110001";
        when 1800 => y_in <= "10000111"; x_in <= "10001000"; z_correct<="0011100010111000";
        when 1801 => y_in <= "10000111"; x_in <= "10001001"; z_correct<="0011100000111111";
        when 1802 => y_in <= "10000111"; x_in <= "10001010"; z_correct<="0011011111000110";
        when 1803 => y_in <= "10000111"; x_in <= "10001011"; z_correct<="0011011101001101";
        when 1804 => y_in <= "10000111"; x_in <= "10001100"; z_correct<="0011011011010100";
        when 1805 => y_in <= "10000111"; x_in <= "10001101"; z_correct<="0011011001011011";
        when 1806 => y_in <= "10000111"; x_in <= "10001110"; z_correct<="0011010111100010";
        when 1807 => y_in <= "10000111"; x_in <= "10001111"; z_correct<="0011010101101001";
        when 1808 => y_in <= "10000111"; x_in <= "10010000"; z_correct<="0011010011110000";
        when 1809 => y_in <= "10000111"; x_in <= "10010001"; z_correct<="0011010001110111";
        when 1810 => y_in <= "10000111"; x_in <= "10010010"; z_correct<="0011001111111110";
        when 1811 => y_in <= "10000111"; x_in <= "10010011"; z_correct<="0011001110000101";
        when 1812 => y_in <= "10000111"; x_in <= "10010100"; z_correct<="0011001100001100";
        when 1813 => y_in <= "10000111"; x_in <= "10010101"; z_correct<="0011001010010011";
        when 1814 => y_in <= "10000111"; x_in <= "10010110"; z_correct<="0011001000011010";
        when 1815 => y_in <= "10000111"; x_in <= "10010111"; z_correct<="0011000110100001";
        when 1816 => y_in <= "10000111"; x_in <= "10011000"; z_correct<="0011000100101000";
        when 1817 => y_in <= "10000111"; x_in <= "10011001"; z_correct<="0011000010101111";
        when 1818 => y_in <= "10000111"; x_in <= "10011010"; z_correct<="0011000000110110";
        when 1819 => y_in <= "10000111"; x_in <= "10011011"; z_correct<="0010111110111101";
        when 1820 => y_in <= "10000111"; x_in <= "10011100"; z_correct<="0010111101000100";
        when 1821 => y_in <= "10000111"; x_in <= "10011101"; z_correct<="0010111011001011";
        when 1822 => y_in <= "10000111"; x_in <= "10011110"; z_correct<="0010111001010010";
        when 1823 => y_in <= "10000111"; x_in <= "10011111"; z_correct<="0010110111011001";
        when 1824 => y_in <= "10000111"; x_in <= "10100000"; z_correct<="0010110101100000";
        when 1825 => y_in <= "10000111"; x_in <= "10100001"; z_correct<="0010110011100111";
        when 1826 => y_in <= "10000111"; x_in <= "10100010"; z_correct<="0010110001101110";
        when 1827 => y_in <= "10000111"; x_in <= "10100011"; z_correct<="0010101111110101";
        when 1828 => y_in <= "10000111"; x_in <= "10100100"; z_correct<="0010101101111100";
        when 1829 => y_in <= "10000111"; x_in <= "10100101"; z_correct<="0010101100000011";
        when 1830 => y_in <= "10000111"; x_in <= "10100110"; z_correct<="0010101010001010";
        when 1831 => y_in <= "10000111"; x_in <= "10100111"; z_correct<="0010101000010001";
        when 1832 => y_in <= "10000111"; x_in <= "10101000"; z_correct<="0010100110011000";
        when 1833 => y_in <= "10000111"; x_in <= "10101001"; z_correct<="0010100100011111";
        when 1834 => y_in <= "10000111"; x_in <= "10101010"; z_correct<="0010100010100110";
        when 1835 => y_in <= "10000111"; x_in <= "10101011"; z_correct<="0010100000101101";
        when 1836 => y_in <= "10000111"; x_in <= "10101100"; z_correct<="0010011110110100";
        when 1837 => y_in <= "10000111"; x_in <= "10101101"; z_correct<="0010011100111011";
        when 1838 => y_in <= "10000111"; x_in <= "10101110"; z_correct<="0010011011000010";
        when 1839 => y_in <= "10000111"; x_in <= "10101111"; z_correct<="0010011001001001";
        when 1840 => y_in <= "10000111"; x_in <= "10110000"; z_correct<="0010010111010000";
        when 1841 => y_in <= "10000111"; x_in <= "10110001"; z_correct<="0010010101010111";
        when 1842 => y_in <= "10000111"; x_in <= "10110010"; z_correct<="0010010011011110";
        when 1843 => y_in <= "10000111"; x_in <= "10110011"; z_correct<="0010010001100101";
        when 1844 => y_in <= "10000111"; x_in <= "10110100"; z_correct<="0010001111101100";
        when 1845 => y_in <= "10000111"; x_in <= "10110101"; z_correct<="0010001101110011";
        when 1846 => y_in <= "10000111"; x_in <= "10110110"; z_correct<="0010001011111010";
        when 1847 => y_in <= "10000111"; x_in <= "10110111"; z_correct<="0010001010000001";
        when 1848 => y_in <= "10000111"; x_in <= "10111000"; z_correct<="0010001000001000";
        when 1849 => y_in <= "10000111"; x_in <= "10111001"; z_correct<="0010000110001111";
        when 1850 => y_in <= "10000111"; x_in <= "10111010"; z_correct<="0010000100010110";
        when 1851 => y_in <= "10000111"; x_in <= "10111011"; z_correct<="0010000010011101";
        when 1852 => y_in <= "10000111"; x_in <= "10111100"; z_correct<="0010000000100100";
        when 1853 => y_in <= "10000111"; x_in <= "10111101"; z_correct<="0001111110101011";
        when 1854 => y_in <= "10000111"; x_in <= "10111110"; z_correct<="0001111100110010";
        when 1855 => y_in <= "10000111"; x_in <= "10111111"; z_correct<="0001111010111001";
        when 1856 => y_in <= "10000111"; x_in <= "11000000"; z_correct<="0001111001000000";
        when 1857 => y_in <= "10000111"; x_in <= "11000001"; z_correct<="0001110111000111";
        when 1858 => y_in <= "10000111"; x_in <= "11000010"; z_correct<="0001110101001110";
        when 1859 => y_in <= "10000111"; x_in <= "11000011"; z_correct<="0001110011010101";
        when 1860 => y_in <= "10000111"; x_in <= "11000100"; z_correct<="0001110001011100";
        when 1861 => y_in <= "10000111"; x_in <= "11000101"; z_correct<="0001101111100011";
        when 1862 => y_in <= "10000111"; x_in <= "11000110"; z_correct<="0001101101101010";
        when 1863 => y_in <= "10000111"; x_in <= "11000111"; z_correct<="0001101011110001";
        when 1864 => y_in <= "10000111"; x_in <= "11001000"; z_correct<="0001101001111000";
        when 1865 => y_in <= "10000111"; x_in <= "11001001"; z_correct<="0001100111111111";
        when 1866 => y_in <= "10000111"; x_in <= "11001010"; z_correct<="0001100110000110";
        when 1867 => y_in <= "10000111"; x_in <= "11001011"; z_correct<="0001100100001101";
        when 1868 => y_in <= "10000111"; x_in <= "11001100"; z_correct<="0001100010010100";
        when 1869 => y_in <= "10000111"; x_in <= "11001101"; z_correct<="0001100000011011";
        when 1870 => y_in <= "10000111"; x_in <= "11001110"; z_correct<="0001011110100010";
        when 1871 => y_in <= "10000111"; x_in <= "11001111"; z_correct<="0001011100101001";
        when 1872 => y_in <= "10000111"; x_in <= "11010000"; z_correct<="0001011010110000";
        when 1873 => y_in <= "10000111"; x_in <= "11010001"; z_correct<="0001011000110111";
        when 1874 => y_in <= "10000111"; x_in <= "11010010"; z_correct<="0001010110111110";
        when 1875 => y_in <= "10000111"; x_in <= "11010011"; z_correct<="0001010101000101";
        when 1876 => y_in <= "10000111"; x_in <= "11010100"; z_correct<="0001010011001100";
        when 1877 => y_in <= "10000111"; x_in <= "11010101"; z_correct<="0001010001010011";
        when 1878 => y_in <= "10000111"; x_in <= "11010110"; z_correct<="0001001111011010";
        when 1879 => y_in <= "10000111"; x_in <= "11010111"; z_correct<="0001001101100001";
        when 1880 => y_in <= "10000111"; x_in <= "11011000"; z_correct<="0001001011101000";
        when 1881 => y_in <= "10000111"; x_in <= "11011001"; z_correct<="0001001001101111";
        when 1882 => y_in <= "10000111"; x_in <= "11011010"; z_correct<="0001000111110110";
        when 1883 => y_in <= "10000111"; x_in <= "11011011"; z_correct<="0001000101111101";
        when 1884 => y_in <= "10000111"; x_in <= "11011100"; z_correct<="0001000100000100";
        when 1885 => y_in <= "10000111"; x_in <= "11011101"; z_correct<="0001000010001011";
        when 1886 => y_in <= "10000111"; x_in <= "11011110"; z_correct<="0001000000010010";
        when 1887 => y_in <= "10000111"; x_in <= "11011111"; z_correct<="0000111110011001";
        when 1888 => y_in <= "10000111"; x_in <= "11100000"; z_correct<="0000111100100000";
        when 1889 => y_in <= "10000111"; x_in <= "11100001"; z_correct<="0000111010100111";
        when 1890 => y_in <= "10000111"; x_in <= "11100010"; z_correct<="0000111000101110";
        when 1891 => y_in <= "10000111"; x_in <= "11100011"; z_correct<="0000110110110101";
        when 1892 => y_in <= "10000111"; x_in <= "11100100"; z_correct<="0000110100111100";
        when 1893 => y_in <= "10000111"; x_in <= "11100101"; z_correct<="0000110011000011";
        when 1894 => y_in <= "10000111"; x_in <= "11100110"; z_correct<="0000110001001010";
        when 1895 => y_in <= "10000111"; x_in <= "11100111"; z_correct<="0000101111010001";
        when 1896 => y_in <= "10000111"; x_in <= "11101000"; z_correct<="0000101101011000";
        when 1897 => y_in <= "10000111"; x_in <= "11101001"; z_correct<="0000101011011111";
        when 1898 => y_in <= "10000111"; x_in <= "11101010"; z_correct<="0000101001100110";
        when 1899 => y_in <= "10000111"; x_in <= "11101011"; z_correct<="0000100111101101";
        when 1900 => y_in <= "10000111"; x_in <= "11101100"; z_correct<="0000100101110100";
        when 1901 => y_in <= "10000111"; x_in <= "11101101"; z_correct<="0000100011111011";
        when 1902 => y_in <= "10000111"; x_in <= "11101110"; z_correct<="0000100010000010";
        when 1903 => y_in <= "10000111"; x_in <= "11101111"; z_correct<="0000100000001001";
        when 1904 => y_in <= "10000111"; x_in <= "11110000"; z_correct<="0000011110010000";
        when 1905 => y_in <= "10000111"; x_in <= "11110001"; z_correct<="0000011100010111";
        when 1906 => y_in <= "10000111"; x_in <= "11110010"; z_correct<="0000011010011110";
        when 1907 => y_in <= "10000111"; x_in <= "11110011"; z_correct<="0000011000100101";
        when 1908 => y_in <= "10000111"; x_in <= "11110100"; z_correct<="0000010110101100";
        when 1909 => y_in <= "10000111"; x_in <= "11110101"; z_correct<="0000010100110011";
        when 1910 => y_in <= "10000111"; x_in <= "11110110"; z_correct<="0000010010111010";
        when 1911 => y_in <= "10000111"; x_in <= "11110111"; z_correct<="0000010001000001";
        when 1912 => y_in <= "10000111"; x_in <= "11111000"; z_correct<="0000001111001000";
        when 1913 => y_in <= "10000111"; x_in <= "11111001"; z_correct<="0000001101001111";
        when 1914 => y_in <= "10000111"; x_in <= "11111010"; z_correct<="0000001011010110";
        when 1915 => y_in <= "10000111"; x_in <= "11111011"; z_correct<="0000001001011101";
        when 1916 => y_in <= "10000111"; x_in <= "11111100"; z_correct<="0000000111100100";
        when 1917 => y_in <= "10000111"; x_in <= "11111101"; z_correct<="0000000101101011";
        when 1918 => y_in <= "10000111"; x_in <= "11111110"; z_correct<="0000000011110010";
        when 1919 => y_in <= "10000111"; x_in <= "11111111"; z_correct<="0000000001111001";
        when 1920 => y_in <= "10000111"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 1921 => y_in <= "10000111"; x_in <= "00000001"; z_correct<="1111111110000111";
        when 1922 => y_in <= "10000111"; x_in <= "00000010"; z_correct<="1111111100001110";
        when 1923 => y_in <= "10000111"; x_in <= "00000011"; z_correct<="1111111010010101";
        when 1924 => y_in <= "10000111"; x_in <= "00000100"; z_correct<="1111111000011100";
        when 1925 => y_in <= "10000111"; x_in <= "00000101"; z_correct<="1111110110100011";
        when 1926 => y_in <= "10000111"; x_in <= "00000110"; z_correct<="1111110100101010";
        when 1927 => y_in <= "10000111"; x_in <= "00000111"; z_correct<="1111110010110001";
        when 1928 => y_in <= "10000111"; x_in <= "00001000"; z_correct<="1111110000111000";
        when 1929 => y_in <= "10000111"; x_in <= "00001001"; z_correct<="1111101110111111";
        when 1930 => y_in <= "10000111"; x_in <= "00001010"; z_correct<="1111101101000110";
        when 1931 => y_in <= "10000111"; x_in <= "00001011"; z_correct<="1111101011001101";
        when 1932 => y_in <= "10000111"; x_in <= "00001100"; z_correct<="1111101001010100";
        when 1933 => y_in <= "10000111"; x_in <= "00001101"; z_correct<="1111100111011011";
        when 1934 => y_in <= "10000111"; x_in <= "00001110"; z_correct<="1111100101100010";
        when 1935 => y_in <= "10000111"; x_in <= "00001111"; z_correct<="1111100011101001";
        when 1936 => y_in <= "10000111"; x_in <= "00010000"; z_correct<="1111100001110000";
        when 1937 => y_in <= "10000111"; x_in <= "00010001"; z_correct<="1111011111110111";
        when 1938 => y_in <= "10000111"; x_in <= "00010010"; z_correct<="1111011101111110";
        when 1939 => y_in <= "10000111"; x_in <= "00010011"; z_correct<="1111011100000101";
        when 1940 => y_in <= "10000111"; x_in <= "00010100"; z_correct<="1111011010001100";
        when 1941 => y_in <= "10000111"; x_in <= "00010101"; z_correct<="1111011000010011";
        when 1942 => y_in <= "10000111"; x_in <= "00010110"; z_correct<="1111010110011010";
        when 1943 => y_in <= "10000111"; x_in <= "00010111"; z_correct<="1111010100100001";
        when 1944 => y_in <= "10000111"; x_in <= "00011000"; z_correct<="1111010010101000";
        when 1945 => y_in <= "10000111"; x_in <= "00011001"; z_correct<="1111010000101111";
        when 1946 => y_in <= "10000111"; x_in <= "00011010"; z_correct<="1111001110110110";
        when 1947 => y_in <= "10000111"; x_in <= "00011011"; z_correct<="1111001100111101";
        when 1948 => y_in <= "10000111"; x_in <= "00011100"; z_correct<="1111001011000100";
        when 1949 => y_in <= "10000111"; x_in <= "00011101"; z_correct<="1111001001001011";
        when 1950 => y_in <= "10000111"; x_in <= "00011110"; z_correct<="1111000111010010";
        when 1951 => y_in <= "10000111"; x_in <= "00011111"; z_correct<="1111000101011001";
        when 1952 => y_in <= "10000111"; x_in <= "00100000"; z_correct<="1111000011100000";
        when 1953 => y_in <= "10000111"; x_in <= "00100001"; z_correct<="1111000001100111";
        when 1954 => y_in <= "10000111"; x_in <= "00100010"; z_correct<="1110111111101110";
        when 1955 => y_in <= "10000111"; x_in <= "00100011"; z_correct<="1110111101110101";
        when 1956 => y_in <= "10000111"; x_in <= "00100100"; z_correct<="1110111011111100";
        when 1957 => y_in <= "10000111"; x_in <= "00100101"; z_correct<="1110111010000011";
        when 1958 => y_in <= "10000111"; x_in <= "00100110"; z_correct<="1110111000001010";
        when 1959 => y_in <= "10000111"; x_in <= "00100111"; z_correct<="1110110110010001";
        when 1960 => y_in <= "10000111"; x_in <= "00101000"; z_correct<="1110110100011000";
        when 1961 => y_in <= "10000111"; x_in <= "00101001"; z_correct<="1110110010011111";
        when 1962 => y_in <= "10000111"; x_in <= "00101010"; z_correct<="1110110000100110";
        when 1963 => y_in <= "10000111"; x_in <= "00101011"; z_correct<="1110101110101101";
        when 1964 => y_in <= "10000111"; x_in <= "00101100"; z_correct<="1110101100110100";
        when 1965 => y_in <= "10000111"; x_in <= "00101101"; z_correct<="1110101010111011";
        when 1966 => y_in <= "10000111"; x_in <= "00101110"; z_correct<="1110101001000010";
        when 1967 => y_in <= "10000111"; x_in <= "00101111"; z_correct<="1110100111001001";
        when 1968 => y_in <= "10000111"; x_in <= "00110000"; z_correct<="1110100101010000";
        when 1969 => y_in <= "10000111"; x_in <= "00110001"; z_correct<="1110100011010111";
        when 1970 => y_in <= "10000111"; x_in <= "00110010"; z_correct<="1110100001011110";
        when 1971 => y_in <= "10000111"; x_in <= "00110011"; z_correct<="1110011111100101";
        when 1972 => y_in <= "10000111"; x_in <= "00110100"; z_correct<="1110011101101100";
        when 1973 => y_in <= "10000111"; x_in <= "00110101"; z_correct<="1110011011110011";
        when 1974 => y_in <= "10000111"; x_in <= "00110110"; z_correct<="1110011001111010";
        when 1975 => y_in <= "10000111"; x_in <= "00110111"; z_correct<="1110011000000001";
        when 1976 => y_in <= "10000111"; x_in <= "00111000"; z_correct<="1110010110001000";
        when 1977 => y_in <= "10000111"; x_in <= "00111001"; z_correct<="1110010100001111";
        when 1978 => y_in <= "10000111"; x_in <= "00111010"; z_correct<="1110010010010110";
        when 1979 => y_in <= "10000111"; x_in <= "00111011"; z_correct<="1110010000011101";
        when 1980 => y_in <= "10000111"; x_in <= "00111100"; z_correct<="1110001110100100";
        when 1981 => y_in <= "10000111"; x_in <= "00111101"; z_correct<="1110001100101011";
        when 1982 => y_in <= "10000111"; x_in <= "00111110"; z_correct<="1110001010110010";
        when 1983 => y_in <= "10000111"; x_in <= "00111111"; z_correct<="1110001000111001";
        when 1984 => y_in <= "10000111"; x_in <= "01000000"; z_correct<="1110000111000000";
        when 1985 => y_in <= "10000111"; x_in <= "01000001"; z_correct<="1110000101000111";
        when 1986 => y_in <= "10000111"; x_in <= "01000010"; z_correct<="1110000011001110";
        when 1987 => y_in <= "10000111"; x_in <= "01000011"; z_correct<="1110000001010101";
        when 1988 => y_in <= "10000111"; x_in <= "01000100"; z_correct<="1101111111011100";
        when 1989 => y_in <= "10000111"; x_in <= "01000101"; z_correct<="1101111101100011";
        when 1990 => y_in <= "10000111"; x_in <= "01000110"; z_correct<="1101111011101010";
        when 1991 => y_in <= "10000111"; x_in <= "01000111"; z_correct<="1101111001110001";
        when 1992 => y_in <= "10000111"; x_in <= "01001000"; z_correct<="1101110111111000";
        when 1993 => y_in <= "10000111"; x_in <= "01001001"; z_correct<="1101110101111111";
        when 1994 => y_in <= "10000111"; x_in <= "01001010"; z_correct<="1101110100000110";
        when 1995 => y_in <= "10000111"; x_in <= "01001011"; z_correct<="1101110010001101";
        when 1996 => y_in <= "10000111"; x_in <= "01001100"; z_correct<="1101110000010100";
        when 1997 => y_in <= "10000111"; x_in <= "01001101"; z_correct<="1101101110011011";
        when 1998 => y_in <= "10000111"; x_in <= "01001110"; z_correct<="1101101100100010";
        when 1999 => y_in <= "10000111"; x_in <= "01001111"; z_correct<="1101101010101001";
        when 2000 => y_in <= "10000111"; x_in <= "01010000"; z_correct<="1101101000110000";
        when 2001 => y_in <= "10000111"; x_in <= "01010001"; z_correct<="1101100110110111";
        when 2002 => y_in <= "10000111"; x_in <= "01010010"; z_correct<="1101100100111110";
        when 2003 => y_in <= "10000111"; x_in <= "01010011"; z_correct<="1101100011000101";
        when 2004 => y_in <= "10000111"; x_in <= "01010100"; z_correct<="1101100001001100";
        when 2005 => y_in <= "10000111"; x_in <= "01010101"; z_correct<="1101011111010011";
        when 2006 => y_in <= "10000111"; x_in <= "01010110"; z_correct<="1101011101011010";
        when 2007 => y_in <= "10000111"; x_in <= "01010111"; z_correct<="1101011011100001";
        when 2008 => y_in <= "10000111"; x_in <= "01011000"; z_correct<="1101011001101000";
        when 2009 => y_in <= "10000111"; x_in <= "01011001"; z_correct<="1101010111101111";
        when 2010 => y_in <= "10000111"; x_in <= "01011010"; z_correct<="1101010101110110";
        when 2011 => y_in <= "10000111"; x_in <= "01011011"; z_correct<="1101010011111101";
        when 2012 => y_in <= "10000111"; x_in <= "01011100"; z_correct<="1101010010000100";
        when 2013 => y_in <= "10000111"; x_in <= "01011101"; z_correct<="1101010000001011";
        when 2014 => y_in <= "10000111"; x_in <= "01011110"; z_correct<="1101001110010010";
        when 2015 => y_in <= "10000111"; x_in <= "01011111"; z_correct<="1101001100011001";
        when 2016 => y_in <= "10000111"; x_in <= "01100000"; z_correct<="1101001010100000";
        when 2017 => y_in <= "10000111"; x_in <= "01100001"; z_correct<="1101001000100111";
        when 2018 => y_in <= "10000111"; x_in <= "01100010"; z_correct<="1101000110101110";
        when 2019 => y_in <= "10000111"; x_in <= "01100011"; z_correct<="1101000100110101";
        when 2020 => y_in <= "10000111"; x_in <= "01100100"; z_correct<="1101000010111100";
        when 2021 => y_in <= "10000111"; x_in <= "01100101"; z_correct<="1101000001000011";
        when 2022 => y_in <= "10000111"; x_in <= "01100110"; z_correct<="1100111111001010";
        when 2023 => y_in <= "10000111"; x_in <= "01100111"; z_correct<="1100111101010001";
        when 2024 => y_in <= "10000111"; x_in <= "01101000"; z_correct<="1100111011011000";
        when 2025 => y_in <= "10000111"; x_in <= "01101001"; z_correct<="1100111001011111";
        when 2026 => y_in <= "10000111"; x_in <= "01101010"; z_correct<="1100110111100110";
        when 2027 => y_in <= "10000111"; x_in <= "01101011"; z_correct<="1100110101101101";
        when 2028 => y_in <= "10000111"; x_in <= "01101100"; z_correct<="1100110011110100";
        when 2029 => y_in <= "10000111"; x_in <= "01101101"; z_correct<="1100110001111011";
        when 2030 => y_in <= "10000111"; x_in <= "01101110"; z_correct<="1100110000000010";
        when 2031 => y_in <= "10000111"; x_in <= "01101111"; z_correct<="1100101110001001";
        when 2032 => y_in <= "10000111"; x_in <= "01110000"; z_correct<="1100101100010000";
        when 2033 => y_in <= "10000111"; x_in <= "01110001"; z_correct<="1100101010010111";
        when 2034 => y_in <= "10000111"; x_in <= "01110010"; z_correct<="1100101000011110";
        when 2035 => y_in <= "10000111"; x_in <= "01110011"; z_correct<="1100100110100101";
        when 2036 => y_in <= "10000111"; x_in <= "01110100"; z_correct<="1100100100101100";
        when 2037 => y_in <= "10000111"; x_in <= "01110101"; z_correct<="1100100010110011";
        when 2038 => y_in <= "10000111"; x_in <= "01110110"; z_correct<="1100100000111010";
        when 2039 => y_in <= "10000111"; x_in <= "01110111"; z_correct<="1100011111000001";
        when 2040 => y_in <= "10000111"; x_in <= "01111000"; z_correct<="1100011101001000";
        when 2041 => y_in <= "10000111"; x_in <= "01111001"; z_correct<="1100011011001111";
        when 2042 => y_in <= "10000111"; x_in <= "01111010"; z_correct<="1100011001010110";
        when 2043 => y_in <= "10000111"; x_in <= "01111011"; z_correct<="1100010111011101";
        when 2044 => y_in <= "10000111"; x_in <= "01111100"; z_correct<="1100010101100100";
        when 2045 => y_in <= "10000111"; x_in <= "01111101"; z_correct<="1100010011101011";
        when 2046 => y_in <= "10000111"; x_in <= "01111110"; z_correct<="1100010001110010";
        when 2047 => y_in <= "10000111"; x_in <= "01111111"; z_correct<="1100001111111001";
        when 2048 => y_in <= "10001000"; x_in <= "10000000"; z_correct<="0011110000000000";
        when 2049 => y_in <= "10001000"; x_in <= "10000001"; z_correct<="0011101110001000";
        when 2050 => y_in <= "10001000"; x_in <= "10000010"; z_correct<="0011101100010000";
        when 2051 => y_in <= "10001000"; x_in <= "10000011"; z_correct<="0011101010011000";
        when 2052 => y_in <= "10001000"; x_in <= "10000100"; z_correct<="0011101000100000";
        when 2053 => y_in <= "10001000"; x_in <= "10000101"; z_correct<="0011100110101000";
        when 2054 => y_in <= "10001000"; x_in <= "10000110"; z_correct<="0011100100110000";
        when 2055 => y_in <= "10001000"; x_in <= "10000111"; z_correct<="0011100010111000";
        when 2056 => y_in <= "10001000"; x_in <= "10001000"; z_correct<="0011100001000000";
        when 2057 => y_in <= "10001000"; x_in <= "10001001"; z_correct<="0011011111001000";
        when 2058 => y_in <= "10001000"; x_in <= "10001010"; z_correct<="0011011101010000";
        when 2059 => y_in <= "10001000"; x_in <= "10001011"; z_correct<="0011011011011000";
        when 2060 => y_in <= "10001000"; x_in <= "10001100"; z_correct<="0011011001100000";
        when 2061 => y_in <= "10001000"; x_in <= "10001101"; z_correct<="0011010111101000";
        when 2062 => y_in <= "10001000"; x_in <= "10001110"; z_correct<="0011010101110000";
        when 2063 => y_in <= "10001000"; x_in <= "10001111"; z_correct<="0011010011111000";
        when 2064 => y_in <= "10001000"; x_in <= "10010000"; z_correct<="0011010010000000";
        when 2065 => y_in <= "10001000"; x_in <= "10010001"; z_correct<="0011010000001000";
        when 2066 => y_in <= "10001000"; x_in <= "10010010"; z_correct<="0011001110010000";
        when 2067 => y_in <= "10001000"; x_in <= "10010011"; z_correct<="0011001100011000";
        when 2068 => y_in <= "10001000"; x_in <= "10010100"; z_correct<="0011001010100000";
        when 2069 => y_in <= "10001000"; x_in <= "10010101"; z_correct<="0011001000101000";
        when 2070 => y_in <= "10001000"; x_in <= "10010110"; z_correct<="0011000110110000";
        when 2071 => y_in <= "10001000"; x_in <= "10010111"; z_correct<="0011000100111000";
        when 2072 => y_in <= "10001000"; x_in <= "10011000"; z_correct<="0011000011000000";
        when 2073 => y_in <= "10001000"; x_in <= "10011001"; z_correct<="0011000001001000";
        when 2074 => y_in <= "10001000"; x_in <= "10011010"; z_correct<="0010111111010000";
        when 2075 => y_in <= "10001000"; x_in <= "10011011"; z_correct<="0010111101011000";
        when 2076 => y_in <= "10001000"; x_in <= "10011100"; z_correct<="0010111011100000";
        when 2077 => y_in <= "10001000"; x_in <= "10011101"; z_correct<="0010111001101000";
        when 2078 => y_in <= "10001000"; x_in <= "10011110"; z_correct<="0010110111110000";
        when 2079 => y_in <= "10001000"; x_in <= "10011111"; z_correct<="0010110101111000";
        when 2080 => y_in <= "10001000"; x_in <= "10100000"; z_correct<="0010110100000000";
        when 2081 => y_in <= "10001000"; x_in <= "10100001"; z_correct<="0010110010001000";
        when 2082 => y_in <= "10001000"; x_in <= "10100010"; z_correct<="0010110000010000";
        when 2083 => y_in <= "10001000"; x_in <= "10100011"; z_correct<="0010101110011000";
        when 2084 => y_in <= "10001000"; x_in <= "10100100"; z_correct<="0010101100100000";
        when 2085 => y_in <= "10001000"; x_in <= "10100101"; z_correct<="0010101010101000";
        when 2086 => y_in <= "10001000"; x_in <= "10100110"; z_correct<="0010101000110000";
        when 2087 => y_in <= "10001000"; x_in <= "10100111"; z_correct<="0010100110111000";
        when 2088 => y_in <= "10001000"; x_in <= "10101000"; z_correct<="0010100101000000";
        when 2089 => y_in <= "10001000"; x_in <= "10101001"; z_correct<="0010100011001000";
        when 2090 => y_in <= "10001000"; x_in <= "10101010"; z_correct<="0010100001010000";
        when 2091 => y_in <= "10001000"; x_in <= "10101011"; z_correct<="0010011111011000";
        when 2092 => y_in <= "10001000"; x_in <= "10101100"; z_correct<="0010011101100000";
        when 2093 => y_in <= "10001000"; x_in <= "10101101"; z_correct<="0010011011101000";
        when 2094 => y_in <= "10001000"; x_in <= "10101110"; z_correct<="0010011001110000";
        when 2095 => y_in <= "10001000"; x_in <= "10101111"; z_correct<="0010010111111000";
        when 2096 => y_in <= "10001000"; x_in <= "10110000"; z_correct<="0010010110000000";
        when 2097 => y_in <= "10001000"; x_in <= "10110001"; z_correct<="0010010100001000";
        when 2098 => y_in <= "10001000"; x_in <= "10110010"; z_correct<="0010010010010000";
        when 2099 => y_in <= "10001000"; x_in <= "10110011"; z_correct<="0010010000011000";
        when 2100 => y_in <= "10001000"; x_in <= "10110100"; z_correct<="0010001110100000";
        when 2101 => y_in <= "10001000"; x_in <= "10110101"; z_correct<="0010001100101000";
        when 2102 => y_in <= "10001000"; x_in <= "10110110"; z_correct<="0010001010110000";
        when 2103 => y_in <= "10001000"; x_in <= "10110111"; z_correct<="0010001000111000";
        when 2104 => y_in <= "10001000"; x_in <= "10111000"; z_correct<="0010000111000000";
        when 2105 => y_in <= "10001000"; x_in <= "10111001"; z_correct<="0010000101001000";
        when 2106 => y_in <= "10001000"; x_in <= "10111010"; z_correct<="0010000011010000";
        when 2107 => y_in <= "10001000"; x_in <= "10111011"; z_correct<="0010000001011000";
        when 2108 => y_in <= "10001000"; x_in <= "10111100"; z_correct<="0001111111100000";
        when 2109 => y_in <= "10001000"; x_in <= "10111101"; z_correct<="0001111101101000";
        when 2110 => y_in <= "10001000"; x_in <= "10111110"; z_correct<="0001111011110000";
        when 2111 => y_in <= "10001000"; x_in <= "10111111"; z_correct<="0001111001111000";
        when 2112 => y_in <= "10001000"; x_in <= "11000000"; z_correct<="0001111000000000";
        when 2113 => y_in <= "10001000"; x_in <= "11000001"; z_correct<="0001110110001000";
        when 2114 => y_in <= "10001000"; x_in <= "11000010"; z_correct<="0001110100010000";
        when 2115 => y_in <= "10001000"; x_in <= "11000011"; z_correct<="0001110010011000";
        when 2116 => y_in <= "10001000"; x_in <= "11000100"; z_correct<="0001110000100000";
        when 2117 => y_in <= "10001000"; x_in <= "11000101"; z_correct<="0001101110101000";
        when 2118 => y_in <= "10001000"; x_in <= "11000110"; z_correct<="0001101100110000";
        when 2119 => y_in <= "10001000"; x_in <= "11000111"; z_correct<="0001101010111000";
        when 2120 => y_in <= "10001000"; x_in <= "11001000"; z_correct<="0001101001000000";
        when 2121 => y_in <= "10001000"; x_in <= "11001001"; z_correct<="0001100111001000";
        when 2122 => y_in <= "10001000"; x_in <= "11001010"; z_correct<="0001100101010000";
        when 2123 => y_in <= "10001000"; x_in <= "11001011"; z_correct<="0001100011011000";
        when 2124 => y_in <= "10001000"; x_in <= "11001100"; z_correct<="0001100001100000";
        when 2125 => y_in <= "10001000"; x_in <= "11001101"; z_correct<="0001011111101000";
        when 2126 => y_in <= "10001000"; x_in <= "11001110"; z_correct<="0001011101110000";
        when 2127 => y_in <= "10001000"; x_in <= "11001111"; z_correct<="0001011011111000";
        when 2128 => y_in <= "10001000"; x_in <= "11010000"; z_correct<="0001011010000000";
        when 2129 => y_in <= "10001000"; x_in <= "11010001"; z_correct<="0001011000001000";
        when 2130 => y_in <= "10001000"; x_in <= "11010010"; z_correct<="0001010110010000";
        when 2131 => y_in <= "10001000"; x_in <= "11010011"; z_correct<="0001010100011000";
        when 2132 => y_in <= "10001000"; x_in <= "11010100"; z_correct<="0001010010100000";
        when 2133 => y_in <= "10001000"; x_in <= "11010101"; z_correct<="0001010000101000";
        when 2134 => y_in <= "10001000"; x_in <= "11010110"; z_correct<="0001001110110000";
        when 2135 => y_in <= "10001000"; x_in <= "11010111"; z_correct<="0001001100111000";
        when 2136 => y_in <= "10001000"; x_in <= "11011000"; z_correct<="0001001011000000";
        when 2137 => y_in <= "10001000"; x_in <= "11011001"; z_correct<="0001001001001000";
        when 2138 => y_in <= "10001000"; x_in <= "11011010"; z_correct<="0001000111010000";
        when 2139 => y_in <= "10001000"; x_in <= "11011011"; z_correct<="0001000101011000";
        when 2140 => y_in <= "10001000"; x_in <= "11011100"; z_correct<="0001000011100000";
        when 2141 => y_in <= "10001000"; x_in <= "11011101"; z_correct<="0001000001101000";
        when 2142 => y_in <= "10001000"; x_in <= "11011110"; z_correct<="0000111111110000";
        when 2143 => y_in <= "10001000"; x_in <= "11011111"; z_correct<="0000111101111000";
        when 2144 => y_in <= "10001000"; x_in <= "11100000"; z_correct<="0000111100000000";
        when 2145 => y_in <= "10001000"; x_in <= "11100001"; z_correct<="0000111010001000";
        when 2146 => y_in <= "10001000"; x_in <= "11100010"; z_correct<="0000111000010000";
        when 2147 => y_in <= "10001000"; x_in <= "11100011"; z_correct<="0000110110011000";
        when 2148 => y_in <= "10001000"; x_in <= "11100100"; z_correct<="0000110100100000";
        when 2149 => y_in <= "10001000"; x_in <= "11100101"; z_correct<="0000110010101000";
        when 2150 => y_in <= "10001000"; x_in <= "11100110"; z_correct<="0000110000110000";
        when 2151 => y_in <= "10001000"; x_in <= "11100111"; z_correct<="0000101110111000";
        when 2152 => y_in <= "10001000"; x_in <= "11101000"; z_correct<="0000101101000000";
        when 2153 => y_in <= "10001000"; x_in <= "11101001"; z_correct<="0000101011001000";
        when 2154 => y_in <= "10001000"; x_in <= "11101010"; z_correct<="0000101001010000";
        when 2155 => y_in <= "10001000"; x_in <= "11101011"; z_correct<="0000100111011000";
        when 2156 => y_in <= "10001000"; x_in <= "11101100"; z_correct<="0000100101100000";
        when 2157 => y_in <= "10001000"; x_in <= "11101101"; z_correct<="0000100011101000";
        when 2158 => y_in <= "10001000"; x_in <= "11101110"; z_correct<="0000100001110000";
        when 2159 => y_in <= "10001000"; x_in <= "11101111"; z_correct<="0000011111111000";
        when 2160 => y_in <= "10001000"; x_in <= "11110000"; z_correct<="0000011110000000";
        when 2161 => y_in <= "10001000"; x_in <= "11110001"; z_correct<="0000011100001000";
        when 2162 => y_in <= "10001000"; x_in <= "11110010"; z_correct<="0000011010010000";
        when 2163 => y_in <= "10001000"; x_in <= "11110011"; z_correct<="0000011000011000";
        when 2164 => y_in <= "10001000"; x_in <= "11110100"; z_correct<="0000010110100000";
        when 2165 => y_in <= "10001000"; x_in <= "11110101"; z_correct<="0000010100101000";
        when 2166 => y_in <= "10001000"; x_in <= "11110110"; z_correct<="0000010010110000";
        when 2167 => y_in <= "10001000"; x_in <= "11110111"; z_correct<="0000010000111000";
        when 2168 => y_in <= "10001000"; x_in <= "11111000"; z_correct<="0000001111000000";
        when 2169 => y_in <= "10001000"; x_in <= "11111001"; z_correct<="0000001101001000";
        when 2170 => y_in <= "10001000"; x_in <= "11111010"; z_correct<="0000001011010000";
        when 2171 => y_in <= "10001000"; x_in <= "11111011"; z_correct<="0000001001011000";
        when 2172 => y_in <= "10001000"; x_in <= "11111100"; z_correct<="0000000111100000";
        when 2173 => y_in <= "10001000"; x_in <= "11111101"; z_correct<="0000000101101000";
        when 2174 => y_in <= "10001000"; x_in <= "11111110"; z_correct<="0000000011110000";
        when 2175 => y_in <= "10001000"; x_in <= "11111111"; z_correct<="0000000001111000";
        when 2176 => y_in <= "10001000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 2177 => y_in <= "10001000"; x_in <= "00000001"; z_correct<="1111111110001000";
        when 2178 => y_in <= "10001000"; x_in <= "00000010"; z_correct<="1111111100010000";
        when 2179 => y_in <= "10001000"; x_in <= "00000011"; z_correct<="1111111010011000";
        when 2180 => y_in <= "10001000"; x_in <= "00000100"; z_correct<="1111111000100000";
        when 2181 => y_in <= "10001000"; x_in <= "00000101"; z_correct<="1111110110101000";
        when 2182 => y_in <= "10001000"; x_in <= "00000110"; z_correct<="1111110100110000";
        when 2183 => y_in <= "10001000"; x_in <= "00000111"; z_correct<="1111110010111000";
        when 2184 => y_in <= "10001000"; x_in <= "00001000"; z_correct<="1111110001000000";
        when 2185 => y_in <= "10001000"; x_in <= "00001001"; z_correct<="1111101111001000";
        when 2186 => y_in <= "10001000"; x_in <= "00001010"; z_correct<="1111101101010000";
        when 2187 => y_in <= "10001000"; x_in <= "00001011"; z_correct<="1111101011011000";
        when 2188 => y_in <= "10001000"; x_in <= "00001100"; z_correct<="1111101001100000";
        when 2189 => y_in <= "10001000"; x_in <= "00001101"; z_correct<="1111100111101000";
        when 2190 => y_in <= "10001000"; x_in <= "00001110"; z_correct<="1111100101110000";
        when 2191 => y_in <= "10001000"; x_in <= "00001111"; z_correct<="1111100011111000";
        when 2192 => y_in <= "10001000"; x_in <= "00010000"; z_correct<="1111100010000000";
        when 2193 => y_in <= "10001000"; x_in <= "00010001"; z_correct<="1111100000001000";
        when 2194 => y_in <= "10001000"; x_in <= "00010010"; z_correct<="1111011110010000";
        when 2195 => y_in <= "10001000"; x_in <= "00010011"; z_correct<="1111011100011000";
        when 2196 => y_in <= "10001000"; x_in <= "00010100"; z_correct<="1111011010100000";
        when 2197 => y_in <= "10001000"; x_in <= "00010101"; z_correct<="1111011000101000";
        when 2198 => y_in <= "10001000"; x_in <= "00010110"; z_correct<="1111010110110000";
        when 2199 => y_in <= "10001000"; x_in <= "00010111"; z_correct<="1111010100111000";
        when 2200 => y_in <= "10001000"; x_in <= "00011000"; z_correct<="1111010011000000";
        when 2201 => y_in <= "10001000"; x_in <= "00011001"; z_correct<="1111010001001000";
        when 2202 => y_in <= "10001000"; x_in <= "00011010"; z_correct<="1111001111010000";
        when 2203 => y_in <= "10001000"; x_in <= "00011011"; z_correct<="1111001101011000";
        when 2204 => y_in <= "10001000"; x_in <= "00011100"; z_correct<="1111001011100000";
        when 2205 => y_in <= "10001000"; x_in <= "00011101"; z_correct<="1111001001101000";
        when 2206 => y_in <= "10001000"; x_in <= "00011110"; z_correct<="1111000111110000";
        when 2207 => y_in <= "10001000"; x_in <= "00011111"; z_correct<="1111000101111000";
        when 2208 => y_in <= "10001000"; x_in <= "00100000"; z_correct<="1111000100000000";
        when 2209 => y_in <= "10001000"; x_in <= "00100001"; z_correct<="1111000010001000";
        when 2210 => y_in <= "10001000"; x_in <= "00100010"; z_correct<="1111000000010000";
        when 2211 => y_in <= "10001000"; x_in <= "00100011"; z_correct<="1110111110011000";
        when 2212 => y_in <= "10001000"; x_in <= "00100100"; z_correct<="1110111100100000";
        when 2213 => y_in <= "10001000"; x_in <= "00100101"; z_correct<="1110111010101000";
        when 2214 => y_in <= "10001000"; x_in <= "00100110"; z_correct<="1110111000110000";
        when 2215 => y_in <= "10001000"; x_in <= "00100111"; z_correct<="1110110110111000";
        when 2216 => y_in <= "10001000"; x_in <= "00101000"; z_correct<="1110110101000000";
        when 2217 => y_in <= "10001000"; x_in <= "00101001"; z_correct<="1110110011001000";
        when 2218 => y_in <= "10001000"; x_in <= "00101010"; z_correct<="1110110001010000";
        when 2219 => y_in <= "10001000"; x_in <= "00101011"; z_correct<="1110101111011000";
        when 2220 => y_in <= "10001000"; x_in <= "00101100"; z_correct<="1110101101100000";
        when 2221 => y_in <= "10001000"; x_in <= "00101101"; z_correct<="1110101011101000";
        when 2222 => y_in <= "10001000"; x_in <= "00101110"; z_correct<="1110101001110000";
        when 2223 => y_in <= "10001000"; x_in <= "00101111"; z_correct<="1110100111111000";
        when 2224 => y_in <= "10001000"; x_in <= "00110000"; z_correct<="1110100110000000";
        when 2225 => y_in <= "10001000"; x_in <= "00110001"; z_correct<="1110100100001000";
        when 2226 => y_in <= "10001000"; x_in <= "00110010"; z_correct<="1110100010010000";
        when 2227 => y_in <= "10001000"; x_in <= "00110011"; z_correct<="1110100000011000";
        when 2228 => y_in <= "10001000"; x_in <= "00110100"; z_correct<="1110011110100000";
        when 2229 => y_in <= "10001000"; x_in <= "00110101"; z_correct<="1110011100101000";
        when 2230 => y_in <= "10001000"; x_in <= "00110110"; z_correct<="1110011010110000";
        when 2231 => y_in <= "10001000"; x_in <= "00110111"; z_correct<="1110011000111000";
        when 2232 => y_in <= "10001000"; x_in <= "00111000"; z_correct<="1110010111000000";
        when 2233 => y_in <= "10001000"; x_in <= "00111001"; z_correct<="1110010101001000";
        when 2234 => y_in <= "10001000"; x_in <= "00111010"; z_correct<="1110010011010000";
        when 2235 => y_in <= "10001000"; x_in <= "00111011"; z_correct<="1110010001011000";
        when 2236 => y_in <= "10001000"; x_in <= "00111100"; z_correct<="1110001111100000";
        when 2237 => y_in <= "10001000"; x_in <= "00111101"; z_correct<="1110001101101000";
        when 2238 => y_in <= "10001000"; x_in <= "00111110"; z_correct<="1110001011110000";
        when 2239 => y_in <= "10001000"; x_in <= "00111111"; z_correct<="1110001001111000";
        when 2240 => y_in <= "10001000"; x_in <= "01000000"; z_correct<="1110001000000000";
        when 2241 => y_in <= "10001000"; x_in <= "01000001"; z_correct<="1110000110001000";
        when 2242 => y_in <= "10001000"; x_in <= "01000010"; z_correct<="1110000100010000";
        when 2243 => y_in <= "10001000"; x_in <= "01000011"; z_correct<="1110000010011000";
        when 2244 => y_in <= "10001000"; x_in <= "01000100"; z_correct<="1110000000100000";
        when 2245 => y_in <= "10001000"; x_in <= "01000101"; z_correct<="1101111110101000";
        when 2246 => y_in <= "10001000"; x_in <= "01000110"; z_correct<="1101111100110000";
        when 2247 => y_in <= "10001000"; x_in <= "01000111"; z_correct<="1101111010111000";
        when 2248 => y_in <= "10001000"; x_in <= "01001000"; z_correct<="1101111001000000";
        when 2249 => y_in <= "10001000"; x_in <= "01001001"; z_correct<="1101110111001000";
        when 2250 => y_in <= "10001000"; x_in <= "01001010"; z_correct<="1101110101010000";
        when 2251 => y_in <= "10001000"; x_in <= "01001011"; z_correct<="1101110011011000";
        when 2252 => y_in <= "10001000"; x_in <= "01001100"; z_correct<="1101110001100000";
        when 2253 => y_in <= "10001000"; x_in <= "01001101"; z_correct<="1101101111101000";
        when 2254 => y_in <= "10001000"; x_in <= "01001110"; z_correct<="1101101101110000";
        when 2255 => y_in <= "10001000"; x_in <= "01001111"; z_correct<="1101101011111000";
        when 2256 => y_in <= "10001000"; x_in <= "01010000"; z_correct<="1101101010000000";
        when 2257 => y_in <= "10001000"; x_in <= "01010001"; z_correct<="1101101000001000";
        when 2258 => y_in <= "10001000"; x_in <= "01010010"; z_correct<="1101100110010000";
        when 2259 => y_in <= "10001000"; x_in <= "01010011"; z_correct<="1101100100011000";
        when 2260 => y_in <= "10001000"; x_in <= "01010100"; z_correct<="1101100010100000";
        when 2261 => y_in <= "10001000"; x_in <= "01010101"; z_correct<="1101100000101000";
        when 2262 => y_in <= "10001000"; x_in <= "01010110"; z_correct<="1101011110110000";
        when 2263 => y_in <= "10001000"; x_in <= "01010111"; z_correct<="1101011100111000";
        when 2264 => y_in <= "10001000"; x_in <= "01011000"; z_correct<="1101011011000000";
        when 2265 => y_in <= "10001000"; x_in <= "01011001"; z_correct<="1101011001001000";
        when 2266 => y_in <= "10001000"; x_in <= "01011010"; z_correct<="1101010111010000";
        when 2267 => y_in <= "10001000"; x_in <= "01011011"; z_correct<="1101010101011000";
        when 2268 => y_in <= "10001000"; x_in <= "01011100"; z_correct<="1101010011100000";
        when 2269 => y_in <= "10001000"; x_in <= "01011101"; z_correct<="1101010001101000";
        when 2270 => y_in <= "10001000"; x_in <= "01011110"; z_correct<="1101001111110000";
        when 2271 => y_in <= "10001000"; x_in <= "01011111"; z_correct<="1101001101111000";
        when 2272 => y_in <= "10001000"; x_in <= "01100000"; z_correct<="1101001100000000";
        when 2273 => y_in <= "10001000"; x_in <= "01100001"; z_correct<="1101001010001000";
        when 2274 => y_in <= "10001000"; x_in <= "01100010"; z_correct<="1101001000010000";
        when 2275 => y_in <= "10001000"; x_in <= "01100011"; z_correct<="1101000110011000";
        when 2276 => y_in <= "10001000"; x_in <= "01100100"; z_correct<="1101000100100000";
        when 2277 => y_in <= "10001000"; x_in <= "01100101"; z_correct<="1101000010101000";
        when 2278 => y_in <= "10001000"; x_in <= "01100110"; z_correct<="1101000000110000";
        when 2279 => y_in <= "10001000"; x_in <= "01100111"; z_correct<="1100111110111000";
        when 2280 => y_in <= "10001000"; x_in <= "01101000"; z_correct<="1100111101000000";
        when 2281 => y_in <= "10001000"; x_in <= "01101001"; z_correct<="1100111011001000";
        when 2282 => y_in <= "10001000"; x_in <= "01101010"; z_correct<="1100111001010000";
        when 2283 => y_in <= "10001000"; x_in <= "01101011"; z_correct<="1100110111011000";
        when 2284 => y_in <= "10001000"; x_in <= "01101100"; z_correct<="1100110101100000";
        when 2285 => y_in <= "10001000"; x_in <= "01101101"; z_correct<="1100110011101000";
        when 2286 => y_in <= "10001000"; x_in <= "01101110"; z_correct<="1100110001110000";
        when 2287 => y_in <= "10001000"; x_in <= "01101111"; z_correct<="1100101111111000";
        when 2288 => y_in <= "10001000"; x_in <= "01110000"; z_correct<="1100101110000000";
        when 2289 => y_in <= "10001000"; x_in <= "01110001"; z_correct<="1100101100001000";
        when 2290 => y_in <= "10001000"; x_in <= "01110010"; z_correct<="1100101010010000";
        when 2291 => y_in <= "10001000"; x_in <= "01110011"; z_correct<="1100101000011000";
        when 2292 => y_in <= "10001000"; x_in <= "01110100"; z_correct<="1100100110100000";
        when 2293 => y_in <= "10001000"; x_in <= "01110101"; z_correct<="1100100100101000";
        when 2294 => y_in <= "10001000"; x_in <= "01110110"; z_correct<="1100100010110000";
        when 2295 => y_in <= "10001000"; x_in <= "01110111"; z_correct<="1100100000111000";
        when 2296 => y_in <= "10001000"; x_in <= "01111000"; z_correct<="1100011111000000";
        when 2297 => y_in <= "10001000"; x_in <= "01111001"; z_correct<="1100011101001000";
        when 2298 => y_in <= "10001000"; x_in <= "01111010"; z_correct<="1100011011010000";
        when 2299 => y_in <= "10001000"; x_in <= "01111011"; z_correct<="1100011001011000";
        when 2300 => y_in <= "10001000"; x_in <= "01111100"; z_correct<="1100010111100000";
        when 2301 => y_in <= "10001000"; x_in <= "01111101"; z_correct<="1100010101101000";
        when 2302 => y_in <= "10001000"; x_in <= "01111110"; z_correct<="1100010011110000";
        when 2303 => y_in <= "10001000"; x_in <= "01111111"; z_correct<="1100010001111000";
        when 2304 => y_in <= "10001001"; x_in <= "10000000"; z_correct<="0011101110000000";
        when 2305 => y_in <= "10001001"; x_in <= "10000001"; z_correct<="0011101100001001";
        when 2306 => y_in <= "10001001"; x_in <= "10000010"; z_correct<="0011101010010010";
        when 2307 => y_in <= "10001001"; x_in <= "10000011"; z_correct<="0011101000011011";
        when 2308 => y_in <= "10001001"; x_in <= "10000100"; z_correct<="0011100110100100";
        when 2309 => y_in <= "10001001"; x_in <= "10000101"; z_correct<="0011100100101101";
        when 2310 => y_in <= "10001001"; x_in <= "10000110"; z_correct<="0011100010110110";
        when 2311 => y_in <= "10001001"; x_in <= "10000111"; z_correct<="0011100000111111";
        when 2312 => y_in <= "10001001"; x_in <= "10001000"; z_correct<="0011011111001000";
        when 2313 => y_in <= "10001001"; x_in <= "10001001"; z_correct<="0011011101010001";
        when 2314 => y_in <= "10001001"; x_in <= "10001010"; z_correct<="0011011011011010";
        when 2315 => y_in <= "10001001"; x_in <= "10001011"; z_correct<="0011011001100011";
        when 2316 => y_in <= "10001001"; x_in <= "10001100"; z_correct<="0011010111101100";
        when 2317 => y_in <= "10001001"; x_in <= "10001101"; z_correct<="0011010101110101";
        when 2318 => y_in <= "10001001"; x_in <= "10001110"; z_correct<="0011010011111110";
        when 2319 => y_in <= "10001001"; x_in <= "10001111"; z_correct<="0011010010000111";
        when 2320 => y_in <= "10001001"; x_in <= "10010000"; z_correct<="0011010000010000";
        when 2321 => y_in <= "10001001"; x_in <= "10010001"; z_correct<="0011001110011001";
        when 2322 => y_in <= "10001001"; x_in <= "10010010"; z_correct<="0011001100100010";
        when 2323 => y_in <= "10001001"; x_in <= "10010011"; z_correct<="0011001010101011";
        when 2324 => y_in <= "10001001"; x_in <= "10010100"; z_correct<="0011001000110100";
        when 2325 => y_in <= "10001001"; x_in <= "10010101"; z_correct<="0011000110111101";
        when 2326 => y_in <= "10001001"; x_in <= "10010110"; z_correct<="0011000101000110";
        when 2327 => y_in <= "10001001"; x_in <= "10010111"; z_correct<="0011000011001111";
        when 2328 => y_in <= "10001001"; x_in <= "10011000"; z_correct<="0011000001011000";
        when 2329 => y_in <= "10001001"; x_in <= "10011001"; z_correct<="0010111111100001";
        when 2330 => y_in <= "10001001"; x_in <= "10011010"; z_correct<="0010111101101010";
        when 2331 => y_in <= "10001001"; x_in <= "10011011"; z_correct<="0010111011110011";
        when 2332 => y_in <= "10001001"; x_in <= "10011100"; z_correct<="0010111001111100";
        when 2333 => y_in <= "10001001"; x_in <= "10011101"; z_correct<="0010111000000101";
        when 2334 => y_in <= "10001001"; x_in <= "10011110"; z_correct<="0010110110001110";
        when 2335 => y_in <= "10001001"; x_in <= "10011111"; z_correct<="0010110100010111";
        when 2336 => y_in <= "10001001"; x_in <= "10100000"; z_correct<="0010110010100000";
        when 2337 => y_in <= "10001001"; x_in <= "10100001"; z_correct<="0010110000101001";
        when 2338 => y_in <= "10001001"; x_in <= "10100010"; z_correct<="0010101110110010";
        when 2339 => y_in <= "10001001"; x_in <= "10100011"; z_correct<="0010101100111011";
        when 2340 => y_in <= "10001001"; x_in <= "10100100"; z_correct<="0010101011000100";
        when 2341 => y_in <= "10001001"; x_in <= "10100101"; z_correct<="0010101001001101";
        when 2342 => y_in <= "10001001"; x_in <= "10100110"; z_correct<="0010100111010110";
        when 2343 => y_in <= "10001001"; x_in <= "10100111"; z_correct<="0010100101011111";
        when 2344 => y_in <= "10001001"; x_in <= "10101000"; z_correct<="0010100011101000";
        when 2345 => y_in <= "10001001"; x_in <= "10101001"; z_correct<="0010100001110001";
        when 2346 => y_in <= "10001001"; x_in <= "10101010"; z_correct<="0010011111111010";
        when 2347 => y_in <= "10001001"; x_in <= "10101011"; z_correct<="0010011110000011";
        when 2348 => y_in <= "10001001"; x_in <= "10101100"; z_correct<="0010011100001100";
        when 2349 => y_in <= "10001001"; x_in <= "10101101"; z_correct<="0010011010010101";
        when 2350 => y_in <= "10001001"; x_in <= "10101110"; z_correct<="0010011000011110";
        when 2351 => y_in <= "10001001"; x_in <= "10101111"; z_correct<="0010010110100111";
        when 2352 => y_in <= "10001001"; x_in <= "10110000"; z_correct<="0010010100110000";
        when 2353 => y_in <= "10001001"; x_in <= "10110001"; z_correct<="0010010010111001";
        when 2354 => y_in <= "10001001"; x_in <= "10110010"; z_correct<="0010010001000010";
        when 2355 => y_in <= "10001001"; x_in <= "10110011"; z_correct<="0010001111001011";
        when 2356 => y_in <= "10001001"; x_in <= "10110100"; z_correct<="0010001101010100";
        when 2357 => y_in <= "10001001"; x_in <= "10110101"; z_correct<="0010001011011101";
        when 2358 => y_in <= "10001001"; x_in <= "10110110"; z_correct<="0010001001100110";
        when 2359 => y_in <= "10001001"; x_in <= "10110111"; z_correct<="0010000111101111";
        when 2360 => y_in <= "10001001"; x_in <= "10111000"; z_correct<="0010000101111000";
        when 2361 => y_in <= "10001001"; x_in <= "10111001"; z_correct<="0010000100000001";
        when 2362 => y_in <= "10001001"; x_in <= "10111010"; z_correct<="0010000010001010";
        when 2363 => y_in <= "10001001"; x_in <= "10111011"; z_correct<="0010000000010011";
        when 2364 => y_in <= "10001001"; x_in <= "10111100"; z_correct<="0001111110011100";
        when 2365 => y_in <= "10001001"; x_in <= "10111101"; z_correct<="0001111100100101";
        when 2366 => y_in <= "10001001"; x_in <= "10111110"; z_correct<="0001111010101110";
        when 2367 => y_in <= "10001001"; x_in <= "10111111"; z_correct<="0001111000110111";
        when 2368 => y_in <= "10001001"; x_in <= "11000000"; z_correct<="0001110111000000";
        when 2369 => y_in <= "10001001"; x_in <= "11000001"; z_correct<="0001110101001001";
        when 2370 => y_in <= "10001001"; x_in <= "11000010"; z_correct<="0001110011010010";
        when 2371 => y_in <= "10001001"; x_in <= "11000011"; z_correct<="0001110001011011";
        when 2372 => y_in <= "10001001"; x_in <= "11000100"; z_correct<="0001101111100100";
        when 2373 => y_in <= "10001001"; x_in <= "11000101"; z_correct<="0001101101101101";
        when 2374 => y_in <= "10001001"; x_in <= "11000110"; z_correct<="0001101011110110";
        when 2375 => y_in <= "10001001"; x_in <= "11000111"; z_correct<="0001101001111111";
        when 2376 => y_in <= "10001001"; x_in <= "11001000"; z_correct<="0001101000001000";
        when 2377 => y_in <= "10001001"; x_in <= "11001001"; z_correct<="0001100110010001";
        when 2378 => y_in <= "10001001"; x_in <= "11001010"; z_correct<="0001100100011010";
        when 2379 => y_in <= "10001001"; x_in <= "11001011"; z_correct<="0001100010100011";
        when 2380 => y_in <= "10001001"; x_in <= "11001100"; z_correct<="0001100000101100";
        when 2381 => y_in <= "10001001"; x_in <= "11001101"; z_correct<="0001011110110101";
        when 2382 => y_in <= "10001001"; x_in <= "11001110"; z_correct<="0001011100111110";
        when 2383 => y_in <= "10001001"; x_in <= "11001111"; z_correct<="0001011011000111";
        when 2384 => y_in <= "10001001"; x_in <= "11010000"; z_correct<="0001011001010000";
        when 2385 => y_in <= "10001001"; x_in <= "11010001"; z_correct<="0001010111011001";
        when 2386 => y_in <= "10001001"; x_in <= "11010010"; z_correct<="0001010101100010";
        when 2387 => y_in <= "10001001"; x_in <= "11010011"; z_correct<="0001010011101011";
        when 2388 => y_in <= "10001001"; x_in <= "11010100"; z_correct<="0001010001110100";
        when 2389 => y_in <= "10001001"; x_in <= "11010101"; z_correct<="0001001111111101";
        when 2390 => y_in <= "10001001"; x_in <= "11010110"; z_correct<="0001001110000110";
        when 2391 => y_in <= "10001001"; x_in <= "11010111"; z_correct<="0001001100001111";
        when 2392 => y_in <= "10001001"; x_in <= "11011000"; z_correct<="0001001010011000";
        when 2393 => y_in <= "10001001"; x_in <= "11011001"; z_correct<="0001001000100001";
        when 2394 => y_in <= "10001001"; x_in <= "11011010"; z_correct<="0001000110101010";
        when 2395 => y_in <= "10001001"; x_in <= "11011011"; z_correct<="0001000100110011";
        when 2396 => y_in <= "10001001"; x_in <= "11011100"; z_correct<="0001000010111100";
        when 2397 => y_in <= "10001001"; x_in <= "11011101"; z_correct<="0001000001000101";
        when 2398 => y_in <= "10001001"; x_in <= "11011110"; z_correct<="0000111111001110";
        when 2399 => y_in <= "10001001"; x_in <= "11011111"; z_correct<="0000111101010111";
        when 2400 => y_in <= "10001001"; x_in <= "11100000"; z_correct<="0000111011100000";
        when 2401 => y_in <= "10001001"; x_in <= "11100001"; z_correct<="0000111001101001";
        when 2402 => y_in <= "10001001"; x_in <= "11100010"; z_correct<="0000110111110010";
        when 2403 => y_in <= "10001001"; x_in <= "11100011"; z_correct<="0000110101111011";
        when 2404 => y_in <= "10001001"; x_in <= "11100100"; z_correct<="0000110100000100";
        when 2405 => y_in <= "10001001"; x_in <= "11100101"; z_correct<="0000110010001101";
        when 2406 => y_in <= "10001001"; x_in <= "11100110"; z_correct<="0000110000010110";
        when 2407 => y_in <= "10001001"; x_in <= "11100111"; z_correct<="0000101110011111";
        when 2408 => y_in <= "10001001"; x_in <= "11101000"; z_correct<="0000101100101000";
        when 2409 => y_in <= "10001001"; x_in <= "11101001"; z_correct<="0000101010110001";
        when 2410 => y_in <= "10001001"; x_in <= "11101010"; z_correct<="0000101000111010";
        when 2411 => y_in <= "10001001"; x_in <= "11101011"; z_correct<="0000100111000011";
        when 2412 => y_in <= "10001001"; x_in <= "11101100"; z_correct<="0000100101001100";
        when 2413 => y_in <= "10001001"; x_in <= "11101101"; z_correct<="0000100011010101";
        when 2414 => y_in <= "10001001"; x_in <= "11101110"; z_correct<="0000100001011110";
        when 2415 => y_in <= "10001001"; x_in <= "11101111"; z_correct<="0000011111100111";
        when 2416 => y_in <= "10001001"; x_in <= "11110000"; z_correct<="0000011101110000";
        when 2417 => y_in <= "10001001"; x_in <= "11110001"; z_correct<="0000011011111001";
        when 2418 => y_in <= "10001001"; x_in <= "11110010"; z_correct<="0000011010000010";
        when 2419 => y_in <= "10001001"; x_in <= "11110011"; z_correct<="0000011000001011";
        when 2420 => y_in <= "10001001"; x_in <= "11110100"; z_correct<="0000010110010100";
        when 2421 => y_in <= "10001001"; x_in <= "11110101"; z_correct<="0000010100011101";
        when 2422 => y_in <= "10001001"; x_in <= "11110110"; z_correct<="0000010010100110";
        when 2423 => y_in <= "10001001"; x_in <= "11110111"; z_correct<="0000010000101111";
        when 2424 => y_in <= "10001001"; x_in <= "11111000"; z_correct<="0000001110111000";
        when 2425 => y_in <= "10001001"; x_in <= "11111001"; z_correct<="0000001101000001";
        when 2426 => y_in <= "10001001"; x_in <= "11111010"; z_correct<="0000001011001010";
        when 2427 => y_in <= "10001001"; x_in <= "11111011"; z_correct<="0000001001010011";
        when 2428 => y_in <= "10001001"; x_in <= "11111100"; z_correct<="0000000111011100";
        when 2429 => y_in <= "10001001"; x_in <= "11111101"; z_correct<="0000000101100101";
        when 2430 => y_in <= "10001001"; x_in <= "11111110"; z_correct<="0000000011101110";
        when 2431 => y_in <= "10001001"; x_in <= "11111111"; z_correct<="0000000001110111";
        when 2432 => y_in <= "10001001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 2433 => y_in <= "10001001"; x_in <= "00000001"; z_correct<="1111111110001001";
        when 2434 => y_in <= "10001001"; x_in <= "00000010"; z_correct<="1111111100010010";
        when 2435 => y_in <= "10001001"; x_in <= "00000011"; z_correct<="1111111010011011";
        when 2436 => y_in <= "10001001"; x_in <= "00000100"; z_correct<="1111111000100100";
        when 2437 => y_in <= "10001001"; x_in <= "00000101"; z_correct<="1111110110101101";
        when 2438 => y_in <= "10001001"; x_in <= "00000110"; z_correct<="1111110100110110";
        when 2439 => y_in <= "10001001"; x_in <= "00000111"; z_correct<="1111110010111111";
        when 2440 => y_in <= "10001001"; x_in <= "00001000"; z_correct<="1111110001001000";
        when 2441 => y_in <= "10001001"; x_in <= "00001001"; z_correct<="1111101111010001";
        when 2442 => y_in <= "10001001"; x_in <= "00001010"; z_correct<="1111101101011010";
        when 2443 => y_in <= "10001001"; x_in <= "00001011"; z_correct<="1111101011100011";
        when 2444 => y_in <= "10001001"; x_in <= "00001100"; z_correct<="1111101001101100";
        when 2445 => y_in <= "10001001"; x_in <= "00001101"; z_correct<="1111100111110101";
        when 2446 => y_in <= "10001001"; x_in <= "00001110"; z_correct<="1111100101111110";
        when 2447 => y_in <= "10001001"; x_in <= "00001111"; z_correct<="1111100100000111";
        when 2448 => y_in <= "10001001"; x_in <= "00010000"; z_correct<="1111100010010000";
        when 2449 => y_in <= "10001001"; x_in <= "00010001"; z_correct<="1111100000011001";
        when 2450 => y_in <= "10001001"; x_in <= "00010010"; z_correct<="1111011110100010";
        when 2451 => y_in <= "10001001"; x_in <= "00010011"; z_correct<="1111011100101011";
        when 2452 => y_in <= "10001001"; x_in <= "00010100"; z_correct<="1111011010110100";
        when 2453 => y_in <= "10001001"; x_in <= "00010101"; z_correct<="1111011000111101";
        when 2454 => y_in <= "10001001"; x_in <= "00010110"; z_correct<="1111010111000110";
        when 2455 => y_in <= "10001001"; x_in <= "00010111"; z_correct<="1111010101001111";
        when 2456 => y_in <= "10001001"; x_in <= "00011000"; z_correct<="1111010011011000";
        when 2457 => y_in <= "10001001"; x_in <= "00011001"; z_correct<="1111010001100001";
        when 2458 => y_in <= "10001001"; x_in <= "00011010"; z_correct<="1111001111101010";
        when 2459 => y_in <= "10001001"; x_in <= "00011011"; z_correct<="1111001101110011";
        when 2460 => y_in <= "10001001"; x_in <= "00011100"; z_correct<="1111001011111100";
        when 2461 => y_in <= "10001001"; x_in <= "00011101"; z_correct<="1111001010000101";
        when 2462 => y_in <= "10001001"; x_in <= "00011110"; z_correct<="1111001000001110";
        when 2463 => y_in <= "10001001"; x_in <= "00011111"; z_correct<="1111000110010111";
        when 2464 => y_in <= "10001001"; x_in <= "00100000"; z_correct<="1111000100100000";
        when 2465 => y_in <= "10001001"; x_in <= "00100001"; z_correct<="1111000010101001";
        when 2466 => y_in <= "10001001"; x_in <= "00100010"; z_correct<="1111000000110010";
        when 2467 => y_in <= "10001001"; x_in <= "00100011"; z_correct<="1110111110111011";
        when 2468 => y_in <= "10001001"; x_in <= "00100100"; z_correct<="1110111101000100";
        when 2469 => y_in <= "10001001"; x_in <= "00100101"; z_correct<="1110111011001101";
        when 2470 => y_in <= "10001001"; x_in <= "00100110"; z_correct<="1110111001010110";
        when 2471 => y_in <= "10001001"; x_in <= "00100111"; z_correct<="1110110111011111";
        when 2472 => y_in <= "10001001"; x_in <= "00101000"; z_correct<="1110110101101000";
        when 2473 => y_in <= "10001001"; x_in <= "00101001"; z_correct<="1110110011110001";
        when 2474 => y_in <= "10001001"; x_in <= "00101010"; z_correct<="1110110001111010";
        when 2475 => y_in <= "10001001"; x_in <= "00101011"; z_correct<="1110110000000011";
        when 2476 => y_in <= "10001001"; x_in <= "00101100"; z_correct<="1110101110001100";
        when 2477 => y_in <= "10001001"; x_in <= "00101101"; z_correct<="1110101100010101";
        when 2478 => y_in <= "10001001"; x_in <= "00101110"; z_correct<="1110101010011110";
        when 2479 => y_in <= "10001001"; x_in <= "00101111"; z_correct<="1110101000100111";
        when 2480 => y_in <= "10001001"; x_in <= "00110000"; z_correct<="1110100110110000";
        when 2481 => y_in <= "10001001"; x_in <= "00110001"; z_correct<="1110100100111001";
        when 2482 => y_in <= "10001001"; x_in <= "00110010"; z_correct<="1110100011000010";
        when 2483 => y_in <= "10001001"; x_in <= "00110011"; z_correct<="1110100001001011";
        when 2484 => y_in <= "10001001"; x_in <= "00110100"; z_correct<="1110011111010100";
        when 2485 => y_in <= "10001001"; x_in <= "00110101"; z_correct<="1110011101011101";
        when 2486 => y_in <= "10001001"; x_in <= "00110110"; z_correct<="1110011011100110";
        when 2487 => y_in <= "10001001"; x_in <= "00110111"; z_correct<="1110011001101111";
        when 2488 => y_in <= "10001001"; x_in <= "00111000"; z_correct<="1110010111111000";
        when 2489 => y_in <= "10001001"; x_in <= "00111001"; z_correct<="1110010110000001";
        when 2490 => y_in <= "10001001"; x_in <= "00111010"; z_correct<="1110010100001010";
        when 2491 => y_in <= "10001001"; x_in <= "00111011"; z_correct<="1110010010010011";
        when 2492 => y_in <= "10001001"; x_in <= "00111100"; z_correct<="1110010000011100";
        when 2493 => y_in <= "10001001"; x_in <= "00111101"; z_correct<="1110001110100101";
        when 2494 => y_in <= "10001001"; x_in <= "00111110"; z_correct<="1110001100101110";
        when 2495 => y_in <= "10001001"; x_in <= "00111111"; z_correct<="1110001010110111";
        when 2496 => y_in <= "10001001"; x_in <= "01000000"; z_correct<="1110001001000000";
        when 2497 => y_in <= "10001001"; x_in <= "01000001"; z_correct<="1110000111001001";
        when 2498 => y_in <= "10001001"; x_in <= "01000010"; z_correct<="1110000101010010";
        when 2499 => y_in <= "10001001"; x_in <= "01000011"; z_correct<="1110000011011011";
        when 2500 => y_in <= "10001001"; x_in <= "01000100"; z_correct<="1110000001100100";
        when 2501 => y_in <= "10001001"; x_in <= "01000101"; z_correct<="1101111111101101";
        when 2502 => y_in <= "10001001"; x_in <= "01000110"; z_correct<="1101111101110110";
        when 2503 => y_in <= "10001001"; x_in <= "01000111"; z_correct<="1101111011111111";
        when 2504 => y_in <= "10001001"; x_in <= "01001000"; z_correct<="1101111010001000";
        when 2505 => y_in <= "10001001"; x_in <= "01001001"; z_correct<="1101111000010001";
        when 2506 => y_in <= "10001001"; x_in <= "01001010"; z_correct<="1101110110011010";
        when 2507 => y_in <= "10001001"; x_in <= "01001011"; z_correct<="1101110100100011";
        when 2508 => y_in <= "10001001"; x_in <= "01001100"; z_correct<="1101110010101100";
        when 2509 => y_in <= "10001001"; x_in <= "01001101"; z_correct<="1101110000110101";
        when 2510 => y_in <= "10001001"; x_in <= "01001110"; z_correct<="1101101110111110";
        when 2511 => y_in <= "10001001"; x_in <= "01001111"; z_correct<="1101101101000111";
        when 2512 => y_in <= "10001001"; x_in <= "01010000"; z_correct<="1101101011010000";
        when 2513 => y_in <= "10001001"; x_in <= "01010001"; z_correct<="1101101001011001";
        when 2514 => y_in <= "10001001"; x_in <= "01010010"; z_correct<="1101100111100010";
        when 2515 => y_in <= "10001001"; x_in <= "01010011"; z_correct<="1101100101101011";
        when 2516 => y_in <= "10001001"; x_in <= "01010100"; z_correct<="1101100011110100";
        when 2517 => y_in <= "10001001"; x_in <= "01010101"; z_correct<="1101100001111101";
        when 2518 => y_in <= "10001001"; x_in <= "01010110"; z_correct<="1101100000000110";
        when 2519 => y_in <= "10001001"; x_in <= "01010111"; z_correct<="1101011110001111";
        when 2520 => y_in <= "10001001"; x_in <= "01011000"; z_correct<="1101011100011000";
        when 2521 => y_in <= "10001001"; x_in <= "01011001"; z_correct<="1101011010100001";
        when 2522 => y_in <= "10001001"; x_in <= "01011010"; z_correct<="1101011000101010";
        when 2523 => y_in <= "10001001"; x_in <= "01011011"; z_correct<="1101010110110011";
        when 2524 => y_in <= "10001001"; x_in <= "01011100"; z_correct<="1101010100111100";
        when 2525 => y_in <= "10001001"; x_in <= "01011101"; z_correct<="1101010011000101";
        when 2526 => y_in <= "10001001"; x_in <= "01011110"; z_correct<="1101010001001110";
        when 2527 => y_in <= "10001001"; x_in <= "01011111"; z_correct<="1101001111010111";
        when 2528 => y_in <= "10001001"; x_in <= "01100000"; z_correct<="1101001101100000";
        when 2529 => y_in <= "10001001"; x_in <= "01100001"; z_correct<="1101001011101001";
        when 2530 => y_in <= "10001001"; x_in <= "01100010"; z_correct<="1101001001110010";
        when 2531 => y_in <= "10001001"; x_in <= "01100011"; z_correct<="1101000111111011";
        when 2532 => y_in <= "10001001"; x_in <= "01100100"; z_correct<="1101000110000100";
        when 2533 => y_in <= "10001001"; x_in <= "01100101"; z_correct<="1101000100001101";
        when 2534 => y_in <= "10001001"; x_in <= "01100110"; z_correct<="1101000010010110";
        when 2535 => y_in <= "10001001"; x_in <= "01100111"; z_correct<="1101000000011111";
        when 2536 => y_in <= "10001001"; x_in <= "01101000"; z_correct<="1100111110101000";
        when 2537 => y_in <= "10001001"; x_in <= "01101001"; z_correct<="1100111100110001";
        when 2538 => y_in <= "10001001"; x_in <= "01101010"; z_correct<="1100111010111010";
        when 2539 => y_in <= "10001001"; x_in <= "01101011"; z_correct<="1100111001000011";
        when 2540 => y_in <= "10001001"; x_in <= "01101100"; z_correct<="1100110111001100";
        when 2541 => y_in <= "10001001"; x_in <= "01101101"; z_correct<="1100110101010101";
        when 2542 => y_in <= "10001001"; x_in <= "01101110"; z_correct<="1100110011011110";
        when 2543 => y_in <= "10001001"; x_in <= "01101111"; z_correct<="1100110001100111";
        when 2544 => y_in <= "10001001"; x_in <= "01110000"; z_correct<="1100101111110000";
        when 2545 => y_in <= "10001001"; x_in <= "01110001"; z_correct<="1100101101111001";
        when 2546 => y_in <= "10001001"; x_in <= "01110010"; z_correct<="1100101100000010";
        when 2547 => y_in <= "10001001"; x_in <= "01110011"; z_correct<="1100101010001011";
        when 2548 => y_in <= "10001001"; x_in <= "01110100"; z_correct<="1100101000010100";
        when 2549 => y_in <= "10001001"; x_in <= "01110101"; z_correct<="1100100110011101";
        when 2550 => y_in <= "10001001"; x_in <= "01110110"; z_correct<="1100100100100110";
        when 2551 => y_in <= "10001001"; x_in <= "01110111"; z_correct<="1100100010101111";
        when 2552 => y_in <= "10001001"; x_in <= "01111000"; z_correct<="1100100000111000";
        when 2553 => y_in <= "10001001"; x_in <= "01111001"; z_correct<="1100011111000001";
        when 2554 => y_in <= "10001001"; x_in <= "01111010"; z_correct<="1100011101001010";
        when 2555 => y_in <= "10001001"; x_in <= "01111011"; z_correct<="1100011011010011";
        when 2556 => y_in <= "10001001"; x_in <= "01111100"; z_correct<="1100011001011100";
        when 2557 => y_in <= "10001001"; x_in <= "01111101"; z_correct<="1100010111100101";
        when 2558 => y_in <= "10001001"; x_in <= "01111110"; z_correct<="1100010101101110";
        when 2559 => y_in <= "10001001"; x_in <= "01111111"; z_correct<="1100010011110111";
        when 2560 => y_in <= "10001010"; x_in <= "10000000"; z_correct<="0011101100000000";
        when 2561 => y_in <= "10001010"; x_in <= "10000001"; z_correct<="0011101010001010";
        when 2562 => y_in <= "10001010"; x_in <= "10000010"; z_correct<="0011101000010100";
        when 2563 => y_in <= "10001010"; x_in <= "10000011"; z_correct<="0011100110011110";
        when 2564 => y_in <= "10001010"; x_in <= "10000100"; z_correct<="0011100100101000";
        when 2565 => y_in <= "10001010"; x_in <= "10000101"; z_correct<="0011100010110010";
        when 2566 => y_in <= "10001010"; x_in <= "10000110"; z_correct<="0011100000111100";
        when 2567 => y_in <= "10001010"; x_in <= "10000111"; z_correct<="0011011111000110";
        when 2568 => y_in <= "10001010"; x_in <= "10001000"; z_correct<="0011011101010000";
        when 2569 => y_in <= "10001010"; x_in <= "10001001"; z_correct<="0011011011011010";
        when 2570 => y_in <= "10001010"; x_in <= "10001010"; z_correct<="0011011001100100";
        when 2571 => y_in <= "10001010"; x_in <= "10001011"; z_correct<="0011010111101110";
        when 2572 => y_in <= "10001010"; x_in <= "10001100"; z_correct<="0011010101111000";
        when 2573 => y_in <= "10001010"; x_in <= "10001101"; z_correct<="0011010100000010";
        when 2574 => y_in <= "10001010"; x_in <= "10001110"; z_correct<="0011010010001100";
        when 2575 => y_in <= "10001010"; x_in <= "10001111"; z_correct<="0011010000010110";
        when 2576 => y_in <= "10001010"; x_in <= "10010000"; z_correct<="0011001110100000";
        when 2577 => y_in <= "10001010"; x_in <= "10010001"; z_correct<="0011001100101010";
        when 2578 => y_in <= "10001010"; x_in <= "10010010"; z_correct<="0011001010110100";
        when 2579 => y_in <= "10001010"; x_in <= "10010011"; z_correct<="0011001000111110";
        when 2580 => y_in <= "10001010"; x_in <= "10010100"; z_correct<="0011000111001000";
        when 2581 => y_in <= "10001010"; x_in <= "10010101"; z_correct<="0011000101010010";
        when 2582 => y_in <= "10001010"; x_in <= "10010110"; z_correct<="0011000011011100";
        when 2583 => y_in <= "10001010"; x_in <= "10010111"; z_correct<="0011000001100110";
        when 2584 => y_in <= "10001010"; x_in <= "10011000"; z_correct<="0010111111110000";
        when 2585 => y_in <= "10001010"; x_in <= "10011001"; z_correct<="0010111101111010";
        when 2586 => y_in <= "10001010"; x_in <= "10011010"; z_correct<="0010111100000100";
        when 2587 => y_in <= "10001010"; x_in <= "10011011"; z_correct<="0010111010001110";
        when 2588 => y_in <= "10001010"; x_in <= "10011100"; z_correct<="0010111000011000";
        when 2589 => y_in <= "10001010"; x_in <= "10011101"; z_correct<="0010110110100010";
        when 2590 => y_in <= "10001010"; x_in <= "10011110"; z_correct<="0010110100101100";
        when 2591 => y_in <= "10001010"; x_in <= "10011111"; z_correct<="0010110010110110";
        when 2592 => y_in <= "10001010"; x_in <= "10100000"; z_correct<="0010110001000000";
        when 2593 => y_in <= "10001010"; x_in <= "10100001"; z_correct<="0010101111001010";
        when 2594 => y_in <= "10001010"; x_in <= "10100010"; z_correct<="0010101101010100";
        when 2595 => y_in <= "10001010"; x_in <= "10100011"; z_correct<="0010101011011110";
        when 2596 => y_in <= "10001010"; x_in <= "10100100"; z_correct<="0010101001101000";
        when 2597 => y_in <= "10001010"; x_in <= "10100101"; z_correct<="0010100111110010";
        when 2598 => y_in <= "10001010"; x_in <= "10100110"; z_correct<="0010100101111100";
        when 2599 => y_in <= "10001010"; x_in <= "10100111"; z_correct<="0010100100000110";
        when 2600 => y_in <= "10001010"; x_in <= "10101000"; z_correct<="0010100010010000";
        when 2601 => y_in <= "10001010"; x_in <= "10101001"; z_correct<="0010100000011010";
        when 2602 => y_in <= "10001010"; x_in <= "10101010"; z_correct<="0010011110100100";
        when 2603 => y_in <= "10001010"; x_in <= "10101011"; z_correct<="0010011100101110";
        when 2604 => y_in <= "10001010"; x_in <= "10101100"; z_correct<="0010011010111000";
        when 2605 => y_in <= "10001010"; x_in <= "10101101"; z_correct<="0010011001000010";
        when 2606 => y_in <= "10001010"; x_in <= "10101110"; z_correct<="0010010111001100";
        when 2607 => y_in <= "10001010"; x_in <= "10101111"; z_correct<="0010010101010110";
        when 2608 => y_in <= "10001010"; x_in <= "10110000"; z_correct<="0010010011100000";
        when 2609 => y_in <= "10001010"; x_in <= "10110001"; z_correct<="0010010001101010";
        when 2610 => y_in <= "10001010"; x_in <= "10110010"; z_correct<="0010001111110100";
        when 2611 => y_in <= "10001010"; x_in <= "10110011"; z_correct<="0010001101111110";
        when 2612 => y_in <= "10001010"; x_in <= "10110100"; z_correct<="0010001100001000";
        when 2613 => y_in <= "10001010"; x_in <= "10110101"; z_correct<="0010001010010010";
        when 2614 => y_in <= "10001010"; x_in <= "10110110"; z_correct<="0010001000011100";
        when 2615 => y_in <= "10001010"; x_in <= "10110111"; z_correct<="0010000110100110";
        when 2616 => y_in <= "10001010"; x_in <= "10111000"; z_correct<="0010000100110000";
        when 2617 => y_in <= "10001010"; x_in <= "10111001"; z_correct<="0010000010111010";
        when 2618 => y_in <= "10001010"; x_in <= "10111010"; z_correct<="0010000001000100";
        when 2619 => y_in <= "10001010"; x_in <= "10111011"; z_correct<="0001111111001110";
        when 2620 => y_in <= "10001010"; x_in <= "10111100"; z_correct<="0001111101011000";
        when 2621 => y_in <= "10001010"; x_in <= "10111101"; z_correct<="0001111011100010";
        when 2622 => y_in <= "10001010"; x_in <= "10111110"; z_correct<="0001111001101100";
        when 2623 => y_in <= "10001010"; x_in <= "10111111"; z_correct<="0001110111110110";
        when 2624 => y_in <= "10001010"; x_in <= "11000000"; z_correct<="0001110110000000";
        when 2625 => y_in <= "10001010"; x_in <= "11000001"; z_correct<="0001110100001010";
        when 2626 => y_in <= "10001010"; x_in <= "11000010"; z_correct<="0001110010010100";
        when 2627 => y_in <= "10001010"; x_in <= "11000011"; z_correct<="0001110000011110";
        when 2628 => y_in <= "10001010"; x_in <= "11000100"; z_correct<="0001101110101000";
        when 2629 => y_in <= "10001010"; x_in <= "11000101"; z_correct<="0001101100110010";
        when 2630 => y_in <= "10001010"; x_in <= "11000110"; z_correct<="0001101010111100";
        when 2631 => y_in <= "10001010"; x_in <= "11000111"; z_correct<="0001101001000110";
        when 2632 => y_in <= "10001010"; x_in <= "11001000"; z_correct<="0001100111010000";
        when 2633 => y_in <= "10001010"; x_in <= "11001001"; z_correct<="0001100101011010";
        when 2634 => y_in <= "10001010"; x_in <= "11001010"; z_correct<="0001100011100100";
        when 2635 => y_in <= "10001010"; x_in <= "11001011"; z_correct<="0001100001101110";
        when 2636 => y_in <= "10001010"; x_in <= "11001100"; z_correct<="0001011111111000";
        when 2637 => y_in <= "10001010"; x_in <= "11001101"; z_correct<="0001011110000010";
        when 2638 => y_in <= "10001010"; x_in <= "11001110"; z_correct<="0001011100001100";
        when 2639 => y_in <= "10001010"; x_in <= "11001111"; z_correct<="0001011010010110";
        when 2640 => y_in <= "10001010"; x_in <= "11010000"; z_correct<="0001011000100000";
        when 2641 => y_in <= "10001010"; x_in <= "11010001"; z_correct<="0001010110101010";
        when 2642 => y_in <= "10001010"; x_in <= "11010010"; z_correct<="0001010100110100";
        when 2643 => y_in <= "10001010"; x_in <= "11010011"; z_correct<="0001010010111110";
        when 2644 => y_in <= "10001010"; x_in <= "11010100"; z_correct<="0001010001001000";
        when 2645 => y_in <= "10001010"; x_in <= "11010101"; z_correct<="0001001111010010";
        when 2646 => y_in <= "10001010"; x_in <= "11010110"; z_correct<="0001001101011100";
        when 2647 => y_in <= "10001010"; x_in <= "11010111"; z_correct<="0001001011100110";
        when 2648 => y_in <= "10001010"; x_in <= "11011000"; z_correct<="0001001001110000";
        when 2649 => y_in <= "10001010"; x_in <= "11011001"; z_correct<="0001000111111010";
        when 2650 => y_in <= "10001010"; x_in <= "11011010"; z_correct<="0001000110000100";
        when 2651 => y_in <= "10001010"; x_in <= "11011011"; z_correct<="0001000100001110";
        when 2652 => y_in <= "10001010"; x_in <= "11011100"; z_correct<="0001000010011000";
        when 2653 => y_in <= "10001010"; x_in <= "11011101"; z_correct<="0001000000100010";
        when 2654 => y_in <= "10001010"; x_in <= "11011110"; z_correct<="0000111110101100";
        when 2655 => y_in <= "10001010"; x_in <= "11011111"; z_correct<="0000111100110110";
        when 2656 => y_in <= "10001010"; x_in <= "11100000"; z_correct<="0000111011000000";
        when 2657 => y_in <= "10001010"; x_in <= "11100001"; z_correct<="0000111001001010";
        when 2658 => y_in <= "10001010"; x_in <= "11100010"; z_correct<="0000110111010100";
        when 2659 => y_in <= "10001010"; x_in <= "11100011"; z_correct<="0000110101011110";
        when 2660 => y_in <= "10001010"; x_in <= "11100100"; z_correct<="0000110011101000";
        when 2661 => y_in <= "10001010"; x_in <= "11100101"; z_correct<="0000110001110010";
        when 2662 => y_in <= "10001010"; x_in <= "11100110"; z_correct<="0000101111111100";
        when 2663 => y_in <= "10001010"; x_in <= "11100111"; z_correct<="0000101110000110";
        when 2664 => y_in <= "10001010"; x_in <= "11101000"; z_correct<="0000101100010000";
        when 2665 => y_in <= "10001010"; x_in <= "11101001"; z_correct<="0000101010011010";
        when 2666 => y_in <= "10001010"; x_in <= "11101010"; z_correct<="0000101000100100";
        when 2667 => y_in <= "10001010"; x_in <= "11101011"; z_correct<="0000100110101110";
        when 2668 => y_in <= "10001010"; x_in <= "11101100"; z_correct<="0000100100111000";
        when 2669 => y_in <= "10001010"; x_in <= "11101101"; z_correct<="0000100011000010";
        when 2670 => y_in <= "10001010"; x_in <= "11101110"; z_correct<="0000100001001100";
        when 2671 => y_in <= "10001010"; x_in <= "11101111"; z_correct<="0000011111010110";
        when 2672 => y_in <= "10001010"; x_in <= "11110000"; z_correct<="0000011101100000";
        when 2673 => y_in <= "10001010"; x_in <= "11110001"; z_correct<="0000011011101010";
        when 2674 => y_in <= "10001010"; x_in <= "11110010"; z_correct<="0000011001110100";
        when 2675 => y_in <= "10001010"; x_in <= "11110011"; z_correct<="0000010111111110";
        when 2676 => y_in <= "10001010"; x_in <= "11110100"; z_correct<="0000010110001000";
        when 2677 => y_in <= "10001010"; x_in <= "11110101"; z_correct<="0000010100010010";
        when 2678 => y_in <= "10001010"; x_in <= "11110110"; z_correct<="0000010010011100";
        when 2679 => y_in <= "10001010"; x_in <= "11110111"; z_correct<="0000010000100110";
        when 2680 => y_in <= "10001010"; x_in <= "11111000"; z_correct<="0000001110110000";
        when 2681 => y_in <= "10001010"; x_in <= "11111001"; z_correct<="0000001100111010";
        when 2682 => y_in <= "10001010"; x_in <= "11111010"; z_correct<="0000001011000100";
        when 2683 => y_in <= "10001010"; x_in <= "11111011"; z_correct<="0000001001001110";
        when 2684 => y_in <= "10001010"; x_in <= "11111100"; z_correct<="0000000111011000";
        when 2685 => y_in <= "10001010"; x_in <= "11111101"; z_correct<="0000000101100010";
        when 2686 => y_in <= "10001010"; x_in <= "11111110"; z_correct<="0000000011101100";
        when 2687 => y_in <= "10001010"; x_in <= "11111111"; z_correct<="0000000001110110";
        when 2688 => y_in <= "10001010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 2689 => y_in <= "10001010"; x_in <= "00000001"; z_correct<="1111111110001010";
        when 2690 => y_in <= "10001010"; x_in <= "00000010"; z_correct<="1111111100010100";
        when 2691 => y_in <= "10001010"; x_in <= "00000011"; z_correct<="1111111010011110";
        when 2692 => y_in <= "10001010"; x_in <= "00000100"; z_correct<="1111111000101000";
        when 2693 => y_in <= "10001010"; x_in <= "00000101"; z_correct<="1111110110110010";
        when 2694 => y_in <= "10001010"; x_in <= "00000110"; z_correct<="1111110100111100";
        when 2695 => y_in <= "10001010"; x_in <= "00000111"; z_correct<="1111110011000110";
        when 2696 => y_in <= "10001010"; x_in <= "00001000"; z_correct<="1111110001010000";
        when 2697 => y_in <= "10001010"; x_in <= "00001001"; z_correct<="1111101111011010";
        when 2698 => y_in <= "10001010"; x_in <= "00001010"; z_correct<="1111101101100100";
        when 2699 => y_in <= "10001010"; x_in <= "00001011"; z_correct<="1111101011101110";
        when 2700 => y_in <= "10001010"; x_in <= "00001100"; z_correct<="1111101001111000";
        when 2701 => y_in <= "10001010"; x_in <= "00001101"; z_correct<="1111101000000010";
        when 2702 => y_in <= "10001010"; x_in <= "00001110"; z_correct<="1111100110001100";
        when 2703 => y_in <= "10001010"; x_in <= "00001111"; z_correct<="1111100100010110";
        when 2704 => y_in <= "10001010"; x_in <= "00010000"; z_correct<="1111100010100000";
        when 2705 => y_in <= "10001010"; x_in <= "00010001"; z_correct<="1111100000101010";
        when 2706 => y_in <= "10001010"; x_in <= "00010010"; z_correct<="1111011110110100";
        when 2707 => y_in <= "10001010"; x_in <= "00010011"; z_correct<="1111011100111110";
        when 2708 => y_in <= "10001010"; x_in <= "00010100"; z_correct<="1111011011001000";
        when 2709 => y_in <= "10001010"; x_in <= "00010101"; z_correct<="1111011001010010";
        when 2710 => y_in <= "10001010"; x_in <= "00010110"; z_correct<="1111010111011100";
        when 2711 => y_in <= "10001010"; x_in <= "00010111"; z_correct<="1111010101100110";
        when 2712 => y_in <= "10001010"; x_in <= "00011000"; z_correct<="1111010011110000";
        when 2713 => y_in <= "10001010"; x_in <= "00011001"; z_correct<="1111010001111010";
        when 2714 => y_in <= "10001010"; x_in <= "00011010"; z_correct<="1111010000000100";
        when 2715 => y_in <= "10001010"; x_in <= "00011011"; z_correct<="1111001110001110";
        when 2716 => y_in <= "10001010"; x_in <= "00011100"; z_correct<="1111001100011000";
        when 2717 => y_in <= "10001010"; x_in <= "00011101"; z_correct<="1111001010100010";
        when 2718 => y_in <= "10001010"; x_in <= "00011110"; z_correct<="1111001000101100";
        when 2719 => y_in <= "10001010"; x_in <= "00011111"; z_correct<="1111000110110110";
        when 2720 => y_in <= "10001010"; x_in <= "00100000"; z_correct<="1111000101000000";
        when 2721 => y_in <= "10001010"; x_in <= "00100001"; z_correct<="1111000011001010";
        when 2722 => y_in <= "10001010"; x_in <= "00100010"; z_correct<="1111000001010100";
        when 2723 => y_in <= "10001010"; x_in <= "00100011"; z_correct<="1110111111011110";
        when 2724 => y_in <= "10001010"; x_in <= "00100100"; z_correct<="1110111101101000";
        when 2725 => y_in <= "10001010"; x_in <= "00100101"; z_correct<="1110111011110010";
        when 2726 => y_in <= "10001010"; x_in <= "00100110"; z_correct<="1110111001111100";
        when 2727 => y_in <= "10001010"; x_in <= "00100111"; z_correct<="1110111000000110";
        when 2728 => y_in <= "10001010"; x_in <= "00101000"; z_correct<="1110110110010000";
        when 2729 => y_in <= "10001010"; x_in <= "00101001"; z_correct<="1110110100011010";
        when 2730 => y_in <= "10001010"; x_in <= "00101010"; z_correct<="1110110010100100";
        when 2731 => y_in <= "10001010"; x_in <= "00101011"; z_correct<="1110110000101110";
        when 2732 => y_in <= "10001010"; x_in <= "00101100"; z_correct<="1110101110111000";
        when 2733 => y_in <= "10001010"; x_in <= "00101101"; z_correct<="1110101101000010";
        when 2734 => y_in <= "10001010"; x_in <= "00101110"; z_correct<="1110101011001100";
        when 2735 => y_in <= "10001010"; x_in <= "00101111"; z_correct<="1110101001010110";
        when 2736 => y_in <= "10001010"; x_in <= "00110000"; z_correct<="1110100111100000";
        when 2737 => y_in <= "10001010"; x_in <= "00110001"; z_correct<="1110100101101010";
        when 2738 => y_in <= "10001010"; x_in <= "00110010"; z_correct<="1110100011110100";
        when 2739 => y_in <= "10001010"; x_in <= "00110011"; z_correct<="1110100001111110";
        when 2740 => y_in <= "10001010"; x_in <= "00110100"; z_correct<="1110100000001000";
        when 2741 => y_in <= "10001010"; x_in <= "00110101"; z_correct<="1110011110010010";
        when 2742 => y_in <= "10001010"; x_in <= "00110110"; z_correct<="1110011100011100";
        when 2743 => y_in <= "10001010"; x_in <= "00110111"; z_correct<="1110011010100110";
        when 2744 => y_in <= "10001010"; x_in <= "00111000"; z_correct<="1110011000110000";
        when 2745 => y_in <= "10001010"; x_in <= "00111001"; z_correct<="1110010110111010";
        when 2746 => y_in <= "10001010"; x_in <= "00111010"; z_correct<="1110010101000100";
        when 2747 => y_in <= "10001010"; x_in <= "00111011"; z_correct<="1110010011001110";
        when 2748 => y_in <= "10001010"; x_in <= "00111100"; z_correct<="1110010001011000";
        when 2749 => y_in <= "10001010"; x_in <= "00111101"; z_correct<="1110001111100010";
        when 2750 => y_in <= "10001010"; x_in <= "00111110"; z_correct<="1110001101101100";
        when 2751 => y_in <= "10001010"; x_in <= "00111111"; z_correct<="1110001011110110";
        when 2752 => y_in <= "10001010"; x_in <= "01000000"; z_correct<="1110001010000000";
        when 2753 => y_in <= "10001010"; x_in <= "01000001"; z_correct<="1110001000001010";
        when 2754 => y_in <= "10001010"; x_in <= "01000010"; z_correct<="1110000110010100";
        when 2755 => y_in <= "10001010"; x_in <= "01000011"; z_correct<="1110000100011110";
        when 2756 => y_in <= "10001010"; x_in <= "01000100"; z_correct<="1110000010101000";
        when 2757 => y_in <= "10001010"; x_in <= "01000101"; z_correct<="1110000000110010";
        when 2758 => y_in <= "10001010"; x_in <= "01000110"; z_correct<="1101111110111100";
        when 2759 => y_in <= "10001010"; x_in <= "01000111"; z_correct<="1101111101000110";
        when 2760 => y_in <= "10001010"; x_in <= "01001000"; z_correct<="1101111011010000";
        when 2761 => y_in <= "10001010"; x_in <= "01001001"; z_correct<="1101111001011010";
        when 2762 => y_in <= "10001010"; x_in <= "01001010"; z_correct<="1101110111100100";
        when 2763 => y_in <= "10001010"; x_in <= "01001011"; z_correct<="1101110101101110";
        when 2764 => y_in <= "10001010"; x_in <= "01001100"; z_correct<="1101110011111000";
        when 2765 => y_in <= "10001010"; x_in <= "01001101"; z_correct<="1101110010000010";
        when 2766 => y_in <= "10001010"; x_in <= "01001110"; z_correct<="1101110000001100";
        when 2767 => y_in <= "10001010"; x_in <= "01001111"; z_correct<="1101101110010110";
        when 2768 => y_in <= "10001010"; x_in <= "01010000"; z_correct<="1101101100100000";
        when 2769 => y_in <= "10001010"; x_in <= "01010001"; z_correct<="1101101010101010";
        when 2770 => y_in <= "10001010"; x_in <= "01010010"; z_correct<="1101101000110100";
        when 2771 => y_in <= "10001010"; x_in <= "01010011"; z_correct<="1101100110111110";
        when 2772 => y_in <= "10001010"; x_in <= "01010100"; z_correct<="1101100101001000";
        when 2773 => y_in <= "10001010"; x_in <= "01010101"; z_correct<="1101100011010010";
        when 2774 => y_in <= "10001010"; x_in <= "01010110"; z_correct<="1101100001011100";
        when 2775 => y_in <= "10001010"; x_in <= "01010111"; z_correct<="1101011111100110";
        when 2776 => y_in <= "10001010"; x_in <= "01011000"; z_correct<="1101011101110000";
        when 2777 => y_in <= "10001010"; x_in <= "01011001"; z_correct<="1101011011111010";
        when 2778 => y_in <= "10001010"; x_in <= "01011010"; z_correct<="1101011010000100";
        when 2779 => y_in <= "10001010"; x_in <= "01011011"; z_correct<="1101011000001110";
        when 2780 => y_in <= "10001010"; x_in <= "01011100"; z_correct<="1101010110011000";
        when 2781 => y_in <= "10001010"; x_in <= "01011101"; z_correct<="1101010100100010";
        when 2782 => y_in <= "10001010"; x_in <= "01011110"; z_correct<="1101010010101100";
        when 2783 => y_in <= "10001010"; x_in <= "01011111"; z_correct<="1101010000110110";
        when 2784 => y_in <= "10001010"; x_in <= "01100000"; z_correct<="1101001111000000";
        when 2785 => y_in <= "10001010"; x_in <= "01100001"; z_correct<="1101001101001010";
        when 2786 => y_in <= "10001010"; x_in <= "01100010"; z_correct<="1101001011010100";
        when 2787 => y_in <= "10001010"; x_in <= "01100011"; z_correct<="1101001001011110";
        when 2788 => y_in <= "10001010"; x_in <= "01100100"; z_correct<="1101000111101000";
        when 2789 => y_in <= "10001010"; x_in <= "01100101"; z_correct<="1101000101110010";
        when 2790 => y_in <= "10001010"; x_in <= "01100110"; z_correct<="1101000011111100";
        when 2791 => y_in <= "10001010"; x_in <= "01100111"; z_correct<="1101000010000110";
        when 2792 => y_in <= "10001010"; x_in <= "01101000"; z_correct<="1101000000010000";
        when 2793 => y_in <= "10001010"; x_in <= "01101001"; z_correct<="1100111110011010";
        when 2794 => y_in <= "10001010"; x_in <= "01101010"; z_correct<="1100111100100100";
        when 2795 => y_in <= "10001010"; x_in <= "01101011"; z_correct<="1100111010101110";
        when 2796 => y_in <= "10001010"; x_in <= "01101100"; z_correct<="1100111000111000";
        when 2797 => y_in <= "10001010"; x_in <= "01101101"; z_correct<="1100110111000010";
        when 2798 => y_in <= "10001010"; x_in <= "01101110"; z_correct<="1100110101001100";
        when 2799 => y_in <= "10001010"; x_in <= "01101111"; z_correct<="1100110011010110";
        when 2800 => y_in <= "10001010"; x_in <= "01110000"; z_correct<="1100110001100000";
        when 2801 => y_in <= "10001010"; x_in <= "01110001"; z_correct<="1100101111101010";
        when 2802 => y_in <= "10001010"; x_in <= "01110010"; z_correct<="1100101101110100";
        when 2803 => y_in <= "10001010"; x_in <= "01110011"; z_correct<="1100101011111110";
        when 2804 => y_in <= "10001010"; x_in <= "01110100"; z_correct<="1100101010001000";
        when 2805 => y_in <= "10001010"; x_in <= "01110101"; z_correct<="1100101000010010";
        when 2806 => y_in <= "10001010"; x_in <= "01110110"; z_correct<="1100100110011100";
        when 2807 => y_in <= "10001010"; x_in <= "01110111"; z_correct<="1100100100100110";
        when 2808 => y_in <= "10001010"; x_in <= "01111000"; z_correct<="1100100010110000";
        when 2809 => y_in <= "10001010"; x_in <= "01111001"; z_correct<="1100100000111010";
        when 2810 => y_in <= "10001010"; x_in <= "01111010"; z_correct<="1100011111000100";
        when 2811 => y_in <= "10001010"; x_in <= "01111011"; z_correct<="1100011101001110";
        when 2812 => y_in <= "10001010"; x_in <= "01111100"; z_correct<="1100011011011000";
        when 2813 => y_in <= "10001010"; x_in <= "01111101"; z_correct<="1100011001100010";
        when 2814 => y_in <= "10001010"; x_in <= "01111110"; z_correct<="1100010111101100";
        when 2815 => y_in <= "10001010"; x_in <= "01111111"; z_correct<="1100010101110110";
        when 2816 => y_in <= "10001011"; x_in <= "10000000"; z_correct<="0011101010000000";
        when 2817 => y_in <= "10001011"; x_in <= "10000001"; z_correct<="0011101000001011";
        when 2818 => y_in <= "10001011"; x_in <= "10000010"; z_correct<="0011100110010110";
        when 2819 => y_in <= "10001011"; x_in <= "10000011"; z_correct<="0011100100100001";
        when 2820 => y_in <= "10001011"; x_in <= "10000100"; z_correct<="0011100010101100";
        when 2821 => y_in <= "10001011"; x_in <= "10000101"; z_correct<="0011100000110111";
        when 2822 => y_in <= "10001011"; x_in <= "10000110"; z_correct<="0011011111000010";
        when 2823 => y_in <= "10001011"; x_in <= "10000111"; z_correct<="0011011101001101";
        when 2824 => y_in <= "10001011"; x_in <= "10001000"; z_correct<="0011011011011000";
        when 2825 => y_in <= "10001011"; x_in <= "10001001"; z_correct<="0011011001100011";
        when 2826 => y_in <= "10001011"; x_in <= "10001010"; z_correct<="0011010111101110";
        when 2827 => y_in <= "10001011"; x_in <= "10001011"; z_correct<="0011010101111001";
        when 2828 => y_in <= "10001011"; x_in <= "10001100"; z_correct<="0011010100000100";
        when 2829 => y_in <= "10001011"; x_in <= "10001101"; z_correct<="0011010010001111";
        when 2830 => y_in <= "10001011"; x_in <= "10001110"; z_correct<="0011010000011010";
        when 2831 => y_in <= "10001011"; x_in <= "10001111"; z_correct<="0011001110100101";
        when 2832 => y_in <= "10001011"; x_in <= "10010000"; z_correct<="0011001100110000";
        when 2833 => y_in <= "10001011"; x_in <= "10010001"; z_correct<="0011001010111011";
        when 2834 => y_in <= "10001011"; x_in <= "10010010"; z_correct<="0011001001000110";
        when 2835 => y_in <= "10001011"; x_in <= "10010011"; z_correct<="0011000111010001";
        when 2836 => y_in <= "10001011"; x_in <= "10010100"; z_correct<="0011000101011100";
        when 2837 => y_in <= "10001011"; x_in <= "10010101"; z_correct<="0011000011100111";
        when 2838 => y_in <= "10001011"; x_in <= "10010110"; z_correct<="0011000001110010";
        when 2839 => y_in <= "10001011"; x_in <= "10010111"; z_correct<="0010111111111101";
        when 2840 => y_in <= "10001011"; x_in <= "10011000"; z_correct<="0010111110001000";
        when 2841 => y_in <= "10001011"; x_in <= "10011001"; z_correct<="0010111100010011";
        when 2842 => y_in <= "10001011"; x_in <= "10011010"; z_correct<="0010111010011110";
        when 2843 => y_in <= "10001011"; x_in <= "10011011"; z_correct<="0010111000101001";
        when 2844 => y_in <= "10001011"; x_in <= "10011100"; z_correct<="0010110110110100";
        when 2845 => y_in <= "10001011"; x_in <= "10011101"; z_correct<="0010110100111111";
        when 2846 => y_in <= "10001011"; x_in <= "10011110"; z_correct<="0010110011001010";
        when 2847 => y_in <= "10001011"; x_in <= "10011111"; z_correct<="0010110001010101";
        when 2848 => y_in <= "10001011"; x_in <= "10100000"; z_correct<="0010101111100000";
        when 2849 => y_in <= "10001011"; x_in <= "10100001"; z_correct<="0010101101101011";
        when 2850 => y_in <= "10001011"; x_in <= "10100010"; z_correct<="0010101011110110";
        when 2851 => y_in <= "10001011"; x_in <= "10100011"; z_correct<="0010101010000001";
        when 2852 => y_in <= "10001011"; x_in <= "10100100"; z_correct<="0010101000001100";
        when 2853 => y_in <= "10001011"; x_in <= "10100101"; z_correct<="0010100110010111";
        when 2854 => y_in <= "10001011"; x_in <= "10100110"; z_correct<="0010100100100010";
        when 2855 => y_in <= "10001011"; x_in <= "10100111"; z_correct<="0010100010101101";
        when 2856 => y_in <= "10001011"; x_in <= "10101000"; z_correct<="0010100000111000";
        when 2857 => y_in <= "10001011"; x_in <= "10101001"; z_correct<="0010011111000011";
        when 2858 => y_in <= "10001011"; x_in <= "10101010"; z_correct<="0010011101001110";
        when 2859 => y_in <= "10001011"; x_in <= "10101011"; z_correct<="0010011011011001";
        when 2860 => y_in <= "10001011"; x_in <= "10101100"; z_correct<="0010011001100100";
        when 2861 => y_in <= "10001011"; x_in <= "10101101"; z_correct<="0010010111101111";
        when 2862 => y_in <= "10001011"; x_in <= "10101110"; z_correct<="0010010101111010";
        when 2863 => y_in <= "10001011"; x_in <= "10101111"; z_correct<="0010010100000101";
        when 2864 => y_in <= "10001011"; x_in <= "10110000"; z_correct<="0010010010010000";
        when 2865 => y_in <= "10001011"; x_in <= "10110001"; z_correct<="0010010000011011";
        when 2866 => y_in <= "10001011"; x_in <= "10110010"; z_correct<="0010001110100110";
        when 2867 => y_in <= "10001011"; x_in <= "10110011"; z_correct<="0010001100110001";
        when 2868 => y_in <= "10001011"; x_in <= "10110100"; z_correct<="0010001010111100";
        when 2869 => y_in <= "10001011"; x_in <= "10110101"; z_correct<="0010001001000111";
        when 2870 => y_in <= "10001011"; x_in <= "10110110"; z_correct<="0010000111010010";
        when 2871 => y_in <= "10001011"; x_in <= "10110111"; z_correct<="0010000101011101";
        when 2872 => y_in <= "10001011"; x_in <= "10111000"; z_correct<="0010000011101000";
        when 2873 => y_in <= "10001011"; x_in <= "10111001"; z_correct<="0010000001110011";
        when 2874 => y_in <= "10001011"; x_in <= "10111010"; z_correct<="0001111111111110";
        when 2875 => y_in <= "10001011"; x_in <= "10111011"; z_correct<="0001111110001001";
        when 2876 => y_in <= "10001011"; x_in <= "10111100"; z_correct<="0001111100010100";
        when 2877 => y_in <= "10001011"; x_in <= "10111101"; z_correct<="0001111010011111";
        when 2878 => y_in <= "10001011"; x_in <= "10111110"; z_correct<="0001111000101010";
        when 2879 => y_in <= "10001011"; x_in <= "10111111"; z_correct<="0001110110110101";
        when 2880 => y_in <= "10001011"; x_in <= "11000000"; z_correct<="0001110101000000";
        when 2881 => y_in <= "10001011"; x_in <= "11000001"; z_correct<="0001110011001011";
        when 2882 => y_in <= "10001011"; x_in <= "11000010"; z_correct<="0001110001010110";
        when 2883 => y_in <= "10001011"; x_in <= "11000011"; z_correct<="0001101111100001";
        when 2884 => y_in <= "10001011"; x_in <= "11000100"; z_correct<="0001101101101100";
        when 2885 => y_in <= "10001011"; x_in <= "11000101"; z_correct<="0001101011110111";
        when 2886 => y_in <= "10001011"; x_in <= "11000110"; z_correct<="0001101010000010";
        when 2887 => y_in <= "10001011"; x_in <= "11000111"; z_correct<="0001101000001101";
        when 2888 => y_in <= "10001011"; x_in <= "11001000"; z_correct<="0001100110011000";
        when 2889 => y_in <= "10001011"; x_in <= "11001001"; z_correct<="0001100100100011";
        when 2890 => y_in <= "10001011"; x_in <= "11001010"; z_correct<="0001100010101110";
        when 2891 => y_in <= "10001011"; x_in <= "11001011"; z_correct<="0001100000111001";
        when 2892 => y_in <= "10001011"; x_in <= "11001100"; z_correct<="0001011111000100";
        when 2893 => y_in <= "10001011"; x_in <= "11001101"; z_correct<="0001011101001111";
        when 2894 => y_in <= "10001011"; x_in <= "11001110"; z_correct<="0001011011011010";
        when 2895 => y_in <= "10001011"; x_in <= "11001111"; z_correct<="0001011001100101";
        when 2896 => y_in <= "10001011"; x_in <= "11010000"; z_correct<="0001010111110000";
        when 2897 => y_in <= "10001011"; x_in <= "11010001"; z_correct<="0001010101111011";
        when 2898 => y_in <= "10001011"; x_in <= "11010010"; z_correct<="0001010100000110";
        when 2899 => y_in <= "10001011"; x_in <= "11010011"; z_correct<="0001010010010001";
        when 2900 => y_in <= "10001011"; x_in <= "11010100"; z_correct<="0001010000011100";
        when 2901 => y_in <= "10001011"; x_in <= "11010101"; z_correct<="0001001110100111";
        when 2902 => y_in <= "10001011"; x_in <= "11010110"; z_correct<="0001001100110010";
        when 2903 => y_in <= "10001011"; x_in <= "11010111"; z_correct<="0001001010111101";
        when 2904 => y_in <= "10001011"; x_in <= "11011000"; z_correct<="0001001001001000";
        when 2905 => y_in <= "10001011"; x_in <= "11011001"; z_correct<="0001000111010011";
        when 2906 => y_in <= "10001011"; x_in <= "11011010"; z_correct<="0001000101011110";
        when 2907 => y_in <= "10001011"; x_in <= "11011011"; z_correct<="0001000011101001";
        when 2908 => y_in <= "10001011"; x_in <= "11011100"; z_correct<="0001000001110100";
        when 2909 => y_in <= "10001011"; x_in <= "11011101"; z_correct<="0000111111111111";
        when 2910 => y_in <= "10001011"; x_in <= "11011110"; z_correct<="0000111110001010";
        when 2911 => y_in <= "10001011"; x_in <= "11011111"; z_correct<="0000111100010101";
        when 2912 => y_in <= "10001011"; x_in <= "11100000"; z_correct<="0000111010100000";
        when 2913 => y_in <= "10001011"; x_in <= "11100001"; z_correct<="0000111000101011";
        when 2914 => y_in <= "10001011"; x_in <= "11100010"; z_correct<="0000110110110110";
        when 2915 => y_in <= "10001011"; x_in <= "11100011"; z_correct<="0000110101000001";
        when 2916 => y_in <= "10001011"; x_in <= "11100100"; z_correct<="0000110011001100";
        when 2917 => y_in <= "10001011"; x_in <= "11100101"; z_correct<="0000110001010111";
        when 2918 => y_in <= "10001011"; x_in <= "11100110"; z_correct<="0000101111100010";
        when 2919 => y_in <= "10001011"; x_in <= "11100111"; z_correct<="0000101101101101";
        when 2920 => y_in <= "10001011"; x_in <= "11101000"; z_correct<="0000101011111000";
        when 2921 => y_in <= "10001011"; x_in <= "11101001"; z_correct<="0000101010000011";
        when 2922 => y_in <= "10001011"; x_in <= "11101010"; z_correct<="0000101000001110";
        when 2923 => y_in <= "10001011"; x_in <= "11101011"; z_correct<="0000100110011001";
        when 2924 => y_in <= "10001011"; x_in <= "11101100"; z_correct<="0000100100100100";
        when 2925 => y_in <= "10001011"; x_in <= "11101101"; z_correct<="0000100010101111";
        when 2926 => y_in <= "10001011"; x_in <= "11101110"; z_correct<="0000100000111010";
        when 2927 => y_in <= "10001011"; x_in <= "11101111"; z_correct<="0000011111000101";
        when 2928 => y_in <= "10001011"; x_in <= "11110000"; z_correct<="0000011101010000";
        when 2929 => y_in <= "10001011"; x_in <= "11110001"; z_correct<="0000011011011011";
        when 2930 => y_in <= "10001011"; x_in <= "11110010"; z_correct<="0000011001100110";
        when 2931 => y_in <= "10001011"; x_in <= "11110011"; z_correct<="0000010111110001";
        when 2932 => y_in <= "10001011"; x_in <= "11110100"; z_correct<="0000010101111100";
        when 2933 => y_in <= "10001011"; x_in <= "11110101"; z_correct<="0000010100000111";
        when 2934 => y_in <= "10001011"; x_in <= "11110110"; z_correct<="0000010010010010";
        when 2935 => y_in <= "10001011"; x_in <= "11110111"; z_correct<="0000010000011101";
        when 2936 => y_in <= "10001011"; x_in <= "11111000"; z_correct<="0000001110101000";
        when 2937 => y_in <= "10001011"; x_in <= "11111001"; z_correct<="0000001100110011";
        when 2938 => y_in <= "10001011"; x_in <= "11111010"; z_correct<="0000001010111110";
        when 2939 => y_in <= "10001011"; x_in <= "11111011"; z_correct<="0000001001001001";
        when 2940 => y_in <= "10001011"; x_in <= "11111100"; z_correct<="0000000111010100";
        when 2941 => y_in <= "10001011"; x_in <= "11111101"; z_correct<="0000000101011111";
        when 2942 => y_in <= "10001011"; x_in <= "11111110"; z_correct<="0000000011101010";
        when 2943 => y_in <= "10001011"; x_in <= "11111111"; z_correct<="0000000001110101";
        when 2944 => y_in <= "10001011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 2945 => y_in <= "10001011"; x_in <= "00000001"; z_correct<="1111111110001011";
        when 2946 => y_in <= "10001011"; x_in <= "00000010"; z_correct<="1111111100010110";
        when 2947 => y_in <= "10001011"; x_in <= "00000011"; z_correct<="1111111010100001";
        when 2948 => y_in <= "10001011"; x_in <= "00000100"; z_correct<="1111111000101100";
        when 2949 => y_in <= "10001011"; x_in <= "00000101"; z_correct<="1111110110110111";
        when 2950 => y_in <= "10001011"; x_in <= "00000110"; z_correct<="1111110101000010";
        when 2951 => y_in <= "10001011"; x_in <= "00000111"; z_correct<="1111110011001101";
        when 2952 => y_in <= "10001011"; x_in <= "00001000"; z_correct<="1111110001011000";
        when 2953 => y_in <= "10001011"; x_in <= "00001001"; z_correct<="1111101111100011";
        when 2954 => y_in <= "10001011"; x_in <= "00001010"; z_correct<="1111101101101110";
        when 2955 => y_in <= "10001011"; x_in <= "00001011"; z_correct<="1111101011111001";
        when 2956 => y_in <= "10001011"; x_in <= "00001100"; z_correct<="1111101010000100";
        when 2957 => y_in <= "10001011"; x_in <= "00001101"; z_correct<="1111101000001111";
        when 2958 => y_in <= "10001011"; x_in <= "00001110"; z_correct<="1111100110011010";
        when 2959 => y_in <= "10001011"; x_in <= "00001111"; z_correct<="1111100100100101";
        when 2960 => y_in <= "10001011"; x_in <= "00010000"; z_correct<="1111100010110000";
        when 2961 => y_in <= "10001011"; x_in <= "00010001"; z_correct<="1111100000111011";
        when 2962 => y_in <= "10001011"; x_in <= "00010010"; z_correct<="1111011111000110";
        when 2963 => y_in <= "10001011"; x_in <= "00010011"; z_correct<="1111011101010001";
        when 2964 => y_in <= "10001011"; x_in <= "00010100"; z_correct<="1111011011011100";
        when 2965 => y_in <= "10001011"; x_in <= "00010101"; z_correct<="1111011001100111";
        when 2966 => y_in <= "10001011"; x_in <= "00010110"; z_correct<="1111010111110010";
        when 2967 => y_in <= "10001011"; x_in <= "00010111"; z_correct<="1111010101111101";
        when 2968 => y_in <= "10001011"; x_in <= "00011000"; z_correct<="1111010100001000";
        when 2969 => y_in <= "10001011"; x_in <= "00011001"; z_correct<="1111010010010011";
        when 2970 => y_in <= "10001011"; x_in <= "00011010"; z_correct<="1111010000011110";
        when 2971 => y_in <= "10001011"; x_in <= "00011011"; z_correct<="1111001110101001";
        when 2972 => y_in <= "10001011"; x_in <= "00011100"; z_correct<="1111001100110100";
        when 2973 => y_in <= "10001011"; x_in <= "00011101"; z_correct<="1111001010111111";
        when 2974 => y_in <= "10001011"; x_in <= "00011110"; z_correct<="1111001001001010";
        when 2975 => y_in <= "10001011"; x_in <= "00011111"; z_correct<="1111000111010101";
        when 2976 => y_in <= "10001011"; x_in <= "00100000"; z_correct<="1111000101100000";
        when 2977 => y_in <= "10001011"; x_in <= "00100001"; z_correct<="1111000011101011";
        when 2978 => y_in <= "10001011"; x_in <= "00100010"; z_correct<="1111000001110110";
        when 2979 => y_in <= "10001011"; x_in <= "00100011"; z_correct<="1111000000000001";
        when 2980 => y_in <= "10001011"; x_in <= "00100100"; z_correct<="1110111110001100";
        when 2981 => y_in <= "10001011"; x_in <= "00100101"; z_correct<="1110111100010111";
        when 2982 => y_in <= "10001011"; x_in <= "00100110"; z_correct<="1110111010100010";
        when 2983 => y_in <= "10001011"; x_in <= "00100111"; z_correct<="1110111000101101";
        when 2984 => y_in <= "10001011"; x_in <= "00101000"; z_correct<="1110110110111000";
        when 2985 => y_in <= "10001011"; x_in <= "00101001"; z_correct<="1110110101000011";
        when 2986 => y_in <= "10001011"; x_in <= "00101010"; z_correct<="1110110011001110";
        when 2987 => y_in <= "10001011"; x_in <= "00101011"; z_correct<="1110110001011001";
        when 2988 => y_in <= "10001011"; x_in <= "00101100"; z_correct<="1110101111100100";
        when 2989 => y_in <= "10001011"; x_in <= "00101101"; z_correct<="1110101101101111";
        when 2990 => y_in <= "10001011"; x_in <= "00101110"; z_correct<="1110101011111010";
        when 2991 => y_in <= "10001011"; x_in <= "00101111"; z_correct<="1110101010000101";
        when 2992 => y_in <= "10001011"; x_in <= "00110000"; z_correct<="1110101000010000";
        when 2993 => y_in <= "10001011"; x_in <= "00110001"; z_correct<="1110100110011011";
        when 2994 => y_in <= "10001011"; x_in <= "00110010"; z_correct<="1110100100100110";
        when 2995 => y_in <= "10001011"; x_in <= "00110011"; z_correct<="1110100010110001";
        when 2996 => y_in <= "10001011"; x_in <= "00110100"; z_correct<="1110100000111100";
        when 2997 => y_in <= "10001011"; x_in <= "00110101"; z_correct<="1110011111000111";
        when 2998 => y_in <= "10001011"; x_in <= "00110110"; z_correct<="1110011101010010";
        when 2999 => y_in <= "10001011"; x_in <= "00110111"; z_correct<="1110011011011101";
        when 3000 => y_in <= "10001011"; x_in <= "00111000"; z_correct<="1110011001101000";
        when 3001 => y_in <= "10001011"; x_in <= "00111001"; z_correct<="1110010111110011";
        when 3002 => y_in <= "10001011"; x_in <= "00111010"; z_correct<="1110010101111110";
        when 3003 => y_in <= "10001011"; x_in <= "00111011"; z_correct<="1110010100001001";
        when 3004 => y_in <= "10001011"; x_in <= "00111100"; z_correct<="1110010010010100";
        when 3005 => y_in <= "10001011"; x_in <= "00111101"; z_correct<="1110010000011111";
        when 3006 => y_in <= "10001011"; x_in <= "00111110"; z_correct<="1110001110101010";
        when 3007 => y_in <= "10001011"; x_in <= "00111111"; z_correct<="1110001100110101";
        when 3008 => y_in <= "10001011"; x_in <= "01000000"; z_correct<="1110001011000000";
        when 3009 => y_in <= "10001011"; x_in <= "01000001"; z_correct<="1110001001001011";
        when 3010 => y_in <= "10001011"; x_in <= "01000010"; z_correct<="1110000111010110";
        when 3011 => y_in <= "10001011"; x_in <= "01000011"; z_correct<="1110000101100001";
        when 3012 => y_in <= "10001011"; x_in <= "01000100"; z_correct<="1110000011101100";
        when 3013 => y_in <= "10001011"; x_in <= "01000101"; z_correct<="1110000001110111";
        when 3014 => y_in <= "10001011"; x_in <= "01000110"; z_correct<="1110000000000010";
        when 3015 => y_in <= "10001011"; x_in <= "01000111"; z_correct<="1101111110001101";
        when 3016 => y_in <= "10001011"; x_in <= "01001000"; z_correct<="1101111100011000";
        when 3017 => y_in <= "10001011"; x_in <= "01001001"; z_correct<="1101111010100011";
        when 3018 => y_in <= "10001011"; x_in <= "01001010"; z_correct<="1101111000101110";
        when 3019 => y_in <= "10001011"; x_in <= "01001011"; z_correct<="1101110110111001";
        when 3020 => y_in <= "10001011"; x_in <= "01001100"; z_correct<="1101110101000100";
        when 3021 => y_in <= "10001011"; x_in <= "01001101"; z_correct<="1101110011001111";
        when 3022 => y_in <= "10001011"; x_in <= "01001110"; z_correct<="1101110001011010";
        when 3023 => y_in <= "10001011"; x_in <= "01001111"; z_correct<="1101101111100101";
        when 3024 => y_in <= "10001011"; x_in <= "01010000"; z_correct<="1101101101110000";
        when 3025 => y_in <= "10001011"; x_in <= "01010001"; z_correct<="1101101011111011";
        when 3026 => y_in <= "10001011"; x_in <= "01010010"; z_correct<="1101101010000110";
        when 3027 => y_in <= "10001011"; x_in <= "01010011"; z_correct<="1101101000010001";
        when 3028 => y_in <= "10001011"; x_in <= "01010100"; z_correct<="1101100110011100";
        when 3029 => y_in <= "10001011"; x_in <= "01010101"; z_correct<="1101100100100111";
        when 3030 => y_in <= "10001011"; x_in <= "01010110"; z_correct<="1101100010110010";
        when 3031 => y_in <= "10001011"; x_in <= "01010111"; z_correct<="1101100000111101";
        when 3032 => y_in <= "10001011"; x_in <= "01011000"; z_correct<="1101011111001000";
        when 3033 => y_in <= "10001011"; x_in <= "01011001"; z_correct<="1101011101010011";
        when 3034 => y_in <= "10001011"; x_in <= "01011010"; z_correct<="1101011011011110";
        when 3035 => y_in <= "10001011"; x_in <= "01011011"; z_correct<="1101011001101001";
        when 3036 => y_in <= "10001011"; x_in <= "01011100"; z_correct<="1101010111110100";
        when 3037 => y_in <= "10001011"; x_in <= "01011101"; z_correct<="1101010101111111";
        when 3038 => y_in <= "10001011"; x_in <= "01011110"; z_correct<="1101010100001010";
        when 3039 => y_in <= "10001011"; x_in <= "01011111"; z_correct<="1101010010010101";
        when 3040 => y_in <= "10001011"; x_in <= "01100000"; z_correct<="1101010000100000";
        when 3041 => y_in <= "10001011"; x_in <= "01100001"; z_correct<="1101001110101011";
        when 3042 => y_in <= "10001011"; x_in <= "01100010"; z_correct<="1101001100110110";
        when 3043 => y_in <= "10001011"; x_in <= "01100011"; z_correct<="1101001011000001";
        when 3044 => y_in <= "10001011"; x_in <= "01100100"; z_correct<="1101001001001100";
        when 3045 => y_in <= "10001011"; x_in <= "01100101"; z_correct<="1101000111010111";
        when 3046 => y_in <= "10001011"; x_in <= "01100110"; z_correct<="1101000101100010";
        when 3047 => y_in <= "10001011"; x_in <= "01100111"; z_correct<="1101000011101101";
        when 3048 => y_in <= "10001011"; x_in <= "01101000"; z_correct<="1101000001111000";
        when 3049 => y_in <= "10001011"; x_in <= "01101001"; z_correct<="1101000000000011";
        when 3050 => y_in <= "10001011"; x_in <= "01101010"; z_correct<="1100111110001110";
        when 3051 => y_in <= "10001011"; x_in <= "01101011"; z_correct<="1100111100011001";
        when 3052 => y_in <= "10001011"; x_in <= "01101100"; z_correct<="1100111010100100";
        when 3053 => y_in <= "10001011"; x_in <= "01101101"; z_correct<="1100111000101111";
        when 3054 => y_in <= "10001011"; x_in <= "01101110"; z_correct<="1100110110111010";
        when 3055 => y_in <= "10001011"; x_in <= "01101111"; z_correct<="1100110101000101";
        when 3056 => y_in <= "10001011"; x_in <= "01110000"; z_correct<="1100110011010000";
        when 3057 => y_in <= "10001011"; x_in <= "01110001"; z_correct<="1100110001011011";
        when 3058 => y_in <= "10001011"; x_in <= "01110010"; z_correct<="1100101111100110";
        when 3059 => y_in <= "10001011"; x_in <= "01110011"; z_correct<="1100101101110001";
        when 3060 => y_in <= "10001011"; x_in <= "01110100"; z_correct<="1100101011111100";
        when 3061 => y_in <= "10001011"; x_in <= "01110101"; z_correct<="1100101010000111";
        when 3062 => y_in <= "10001011"; x_in <= "01110110"; z_correct<="1100101000010010";
        when 3063 => y_in <= "10001011"; x_in <= "01110111"; z_correct<="1100100110011101";
        when 3064 => y_in <= "10001011"; x_in <= "01111000"; z_correct<="1100100100101000";
        when 3065 => y_in <= "10001011"; x_in <= "01111001"; z_correct<="1100100010110011";
        when 3066 => y_in <= "10001011"; x_in <= "01111010"; z_correct<="1100100000111110";
        when 3067 => y_in <= "10001011"; x_in <= "01111011"; z_correct<="1100011111001001";
        when 3068 => y_in <= "10001011"; x_in <= "01111100"; z_correct<="1100011101010100";
        when 3069 => y_in <= "10001011"; x_in <= "01111101"; z_correct<="1100011011011111";
        when 3070 => y_in <= "10001011"; x_in <= "01111110"; z_correct<="1100011001101010";
        when 3071 => y_in <= "10001011"; x_in <= "01111111"; z_correct<="1100010111110101";
        when 3072 => y_in <= "10001100"; x_in <= "10000000"; z_correct<="0011101000000000";
        when 3073 => y_in <= "10001100"; x_in <= "10000001"; z_correct<="0011100110001100";
        when 3074 => y_in <= "10001100"; x_in <= "10000010"; z_correct<="0011100100011000";
        when 3075 => y_in <= "10001100"; x_in <= "10000011"; z_correct<="0011100010100100";
        when 3076 => y_in <= "10001100"; x_in <= "10000100"; z_correct<="0011100000110000";
        when 3077 => y_in <= "10001100"; x_in <= "10000101"; z_correct<="0011011110111100";
        when 3078 => y_in <= "10001100"; x_in <= "10000110"; z_correct<="0011011101001000";
        when 3079 => y_in <= "10001100"; x_in <= "10000111"; z_correct<="0011011011010100";
        when 3080 => y_in <= "10001100"; x_in <= "10001000"; z_correct<="0011011001100000";
        when 3081 => y_in <= "10001100"; x_in <= "10001001"; z_correct<="0011010111101100";
        when 3082 => y_in <= "10001100"; x_in <= "10001010"; z_correct<="0011010101111000";
        when 3083 => y_in <= "10001100"; x_in <= "10001011"; z_correct<="0011010100000100";
        when 3084 => y_in <= "10001100"; x_in <= "10001100"; z_correct<="0011010010010000";
        when 3085 => y_in <= "10001100"; x_in <= "10001101"; z_correct<="0011010000011100";
        when 3086 => y_in <= "10001100"; x_in <= "10001110"; z_correct<="0011001110101000";
        when 3087 => y_in <= "10001100"; x_in <= "10001111"; z_correct<="0011001100110100";
        when 3088 => y_in <= "10001100"; x_in <= "10010000"; z_correct<="0011001011000000";
        when 3089 => y_in <= "10001100"; x_in <= "10010001"; z_correct<="0011001001001100";
        when 3090 => y_in <= "10001100"; x_in <= "10010010"; z_correct<="0011000111011000";
        when 3091 => y_in <= "10001100"; x_in <= "10010011"; z_correct<="0011000101100100";
        when 3092 => y_in <= "10001100"; x_in <= "10010100"; z_correct<="0011000011110000";
        when 3093 => y_in <= "10001100"; x_in <= "10010101"; z_correct<="0011000001111100";
        when 3094 => y_in <= "10001100"; x_in <= "10010110"; z_correct<="0011000000001000";
        when 3095 => y_in <= "10001100"; x_in <= "10010111"; z_correct<="0010111110010100";
        when 3096 => y_in <= "10001100"; x_in <= "10011000"; z_correct<="0010111100100000";
        when 3097 => y_in <= "10001100"; x_in <= "10011001"; z_correct<="0010111010101100";
        when 3098 => y_in <= "10001100"; x_in <= "10011010"; z_correct<="0010111000111000";
        when 3099 => y_in <= "10001100"; x_in <= "10011011"; z_correct<="0010110111000100";
        when 3100 => y_in <= "10001100"; x_in <= "10011100"; z_correct<="0010110101010000";
        when 3101 => y_in <= "10001100"; x_in <= "10011101"; z_correct<="0010110011011100";
        when 3102 => y_in <= "10001100"; x_in <= "10011110"; z_correct<="0010110001101000";
        when 3103 => y_in <= "10001100"; x_in <= "10011111"; z_correct<="0010101111110100";
        when 3104 => y_in <= "10001100"; x_in <= "10100000"; z_correct<="0010101110000000";
        when 3105 => y_in <= "10001100"; x_in <= "10100001"; z_correct<="0010101100001100";
        when 3106 => y_in <= "10001100"; x_in <= "10100010"; z_correct<="0010101010011000";
        when 3107 => y_in <= "10001100"; x_in <= "10100011"; z_correct<="0010101000100100";
        when 3108 => y_in <= "10001100"; x_in <= "10100100"; z_correct<="0010100110110000";
        when 3109 => y_in <= "10001100"; x_in <= "10100101"; z_correct<="0010100100111100";
        when 3110 => y_in <= "10001100"; x_in <= "10100110"; z_correct<="0010100011001000";
        when 3111 => y_in <= "10001100"; x_in <= "10100111"; z_correct<="0010100001010100";
        when 3112 => y_in <= "10001100"; x_in <= "10101000"; z_correct<="0010011111100000";
        when 3113 => y_in <= "10001100"; x_in <= "10101001"; z_correct<="0010011101101100";
        when 3114 => y_in <= "10001100"; x_in <= "10101010"; z_correct<="0010011011111000";
        when 3115 => y_in <= "10001100"; x_in <= "10101011"; z_correct<="0010011010000100";
        when 3116 => y_in <= "10001100"; x_in <= "10101100"; z_correct<="0010011000010000";
        when 3117 => y_in <= "10001100"; x_in <= "10101101"; z_correct<="0010010110011100";
        when 3118 => y_in <= "10001100"; x_in <= "10101110"; z_correct<="0010010100101000";
        when 3119 => y_in <= "10001100"; x_in <= "10101111"; z_correct<="0010010010110100";
        when 3120 => y_in <= "10001100"; x_in <= "10110000"; z_correct<="0010010001000000";
        when 3121 => y_in <= "10001100"; x_in <= "10110001"; z_correct<="0010001111001100";
        when 3122 => y_in <= "10001100"; x_in <= "10110010"; z_correct<="0010001101011000";
        when 3123 => y_in <= "10001100"; x_in <= "10110011"; z_correct<="0010001011100100";
        when 3124 => y_in <= "10001100"; x_in <= "10110100"; z_correct<="0010001001110000";
        when 3125 => y_in <= "10001100"; x_in <= "10110101"; z_correct<="0010000111111100";
        when 3126 => y_in <= "10001100"; x_in <= "10110110"; z_correct<="0010000110001000";
        when 3127 => y_in <= "10001100"; x_in <= "10110111"; z_correct<="0010000100010100";
        when 3128 => y_in <= "10001100"; x_in <= "10111000"; z_correct<="0010000010100000";
        when 3129 => y_in <= "10001100"; x_in <= "10111001"; z_correct<="0010000000101100";
        when 3130 => y_in <= "10001100"; x_in <= "10111010"; z_correct<="0001111110111000";
        when 3131 => y_in <= "10001100"; x_in <= "10111011"; z_correct<="0001111101000100";
        when 3132 => y_in <= "10001100"; x_in <= "10111100"; z_correct<="0001111011010000";
        when 3133 => y_in <= "10001100"; x_in <= "10111101"; z_correct<="0001111001011100";
        when 3134 => y_in <= "10001100"; x_in <= "10111110"; z_correct<="0001110111101000";
        when 3135 => y_in <= "10001100"; x_in <= "10111111"; z_correct<="0001110101110100";
        when 3136 => y_in <= "10001100"; x_in <= "11000000"; z_correct<="0001110100000000";
        when 3137 => y_in <= "10001100"; x_in <= "11000001"; z_correct<="0001110010001100";
        when 3138 => y_in <= "10001100"; x_in <= "11000010"; z_correct<="0001110000011000";
        when 3139 => y_in <= "10001100"; x_in <= "11000011"; z_correct<="0001101110100100";
        when 3140 => y_in <= "10001100"; x_in <= "11000100"; z_correct<="0001101100110000";
        when 3141 => y_in <= "10001100"; x_in <= "11000101"; z_correct<="0001101010111100";
        when 3142 => y_in <= "10001100"; x_in <= "11000110"; z_correct<="0001101001001000";
        when 3143 => y_in <= "10001100"; x_in <= "11000111"; z_correct<="0001100111010100";
        when 3144 => y_in <= "10001100"; x_in <= "11001000"; z_correct<="0001100101100000";
        when 3145 => y_in <= "10001100"; x_in <= "11001001"; z_correct<="0001100011101100";
        when 3146 => y_in <= "10001100"; x_in <= "11001010"; z_correct<="0001100001111000";
        when 3147 => y_in <= "10001100"; x_in <= "11001011"; z_correct<="0001100000000100";
        when 3148 => y_in <= "10001100"; x_in <= "11001100"; z_correct<="0001011110010000";
        when 3149 => y_in <= "10001100"; x_in <= "11001101"; z_correct<="0001011100011100";
        when 3150 => y_in <= "10001100"; x_in <= "11001110"; z_correct<="0001011010101000";
        when 3151 => y_in <= "10001100"; x_in <= "11001111"; z_correct<="0001011000110100";
        when 3152 => y_in <= "10001100"; x_in <= "11010000"; z_correct<="0001010111000000";
        when 3153 => y_in <= "10001100"; x_in <= "11010001"; z_correct<="0001010101001100";
        when 3154 => y_in <= "10001100"; x_in <= "11010010"; z_correct<="0001010011011000";
        when 3155 => y_in <= "10001100"; x_in <= "11010011"; z_correct<="0001010001100100";
        when 3156 => y_in <= "10001100"; x_in <= "11010100"; z_correct<="0001001111110000";
        when 3157 => y_in <= "10001100"; x_in <= "11010101"; z_correct<="0001001101111100";
        when 3158 => y_in <= "10001100"; x_in <= "11010110"; z_correct<="0001001100001000";
        when 3159 => y_in <= "10001100"; x_in <= "11010111"; z_correct<="0001001010010100";
        when 3160 => y_in <= "10001100"; x_in <= "11011000"; z_correct<="0001001000100000";
        when 3161 => y_in <= "10001100"; x_in <= "11011001"; z_correct<="0001000110101100";
        when 3162 => y_in <= "10001100"; x_in <= "11011010"; z_correct<="0001000100111000";
        when 3163 => y_in <= "10001100"; x_in <= "11011011"; z_correct<="0001000011000100";
        when 3164 => y_in <= "10001100"; x_in <= "11011100"; z_correct<="0001000001010000";
        when 3165 => y_in <= "10001100"; x_in <= "11011101"; z_correct<="0000111111011100";
        when 3166 => y_in <= "10001100"; x_in <= "11011110"; z_correct<="0000111101101000";
        when 3167 => y_in <= "10001100"; x_in <= "11011111"; z_correct<="0000111011110100";
        when 3168 => y_in <= "10001100"; x_in <= "11100000"; z_correct<="0000111010000000";
        when 3169 => y_in <= "10001100"; x_in <= "11100001"; z_correct<="0000111000001100";
        when 3170 => y_in <= "10001100"; x_in <= "11100010"; z_correct<="0000110110011000";
        when 3171 => y_in <= "10001100"; x_in <= "11100011"; z_correct<="0000110100100100";
        when 3172 => y_in <= "10001100"; x_in <= "11100100"; z_correct<="0000110010110000";
        when 3173 => y_in <= "10001100"; x_in <= "11100101"; z_correct<="0000110000111100";
        when 3174 => y_in <= "10001100"; x_in <= "11100110"; z_correct<="0000101111001000";
        when 3175 => y_in <= "10001100"; x_in <= "11100111"; z_correct<="0000101101010100";
        when 3176 => y_in <= "10001100"; x_in <= "11101000"; z_correct<="0000101011100000";
        when 3177 => y_in <= "10001100"; x_in <= "11101001"; z_correct<="0000101001101100";
        when 3178 => y_in <= "10001100"; x_in <= "11101010"; z_correct<="0000100111111000";
        when 3179 => y_in <= "10001100"; x_in <= "11101011"; z_correct<="0000100110000100";
        when 3180 => y_in <= "10001100"; x_in <= "11101100"; z_correct<="0000100100010000";
        when 3181 => y_in <= "10001100"; x_in <= "11101101"; z_correct<="0000100010011100";
        when 3182 => y_in <= "10001100"; x_in <= "11101110"; z_correct<="0000100000101000";
        when 3183 => y_in <= "10001100"; x_in <= "11101111"; z_correct<="0000011110110100";
        when 3184 => y_in <= "10001100"; x_in <= "11110000"; z_correct<="0000011101000000";
        when 3185 => y_in <= "10001100"; x_in <= "11110001"; z_correct<="0000011011001100";
        when 3186 => y_in <= "10001100"; x_in <= "11110010"; z_correct<="0000011001011000";
        when 3187 => y_in <= "10001100"; x_in <= "11110011"; z_correct<="0000010111100100";
        when 3188 => y_in <= "10001100"; x_in <= "11110100"; z_correct<="0000010101110000";
        when 3189 => y_in <= "10001100"; x_in <= "11110101"; z_correct<="0000010011111100";
        when 3190 => y_in <= "10001100"; x_in <= "11110110"; z_correct<="0000010010001000";
        when 3191 => y_in <= "10001100"; x_in <= "11110111"; z_correct<="0000010000010100";
        when 3192 => y_in <= "10001100"; x_in <= "11111000"; z_correct<="0000001110100000";
        when 3193 => y_in <= "10001100"; x_in <= "11111001"; z_correct<="0000001100101100";
        when 3194 => y_in <= "10001100"; x_in <= "11111010"; z_correct<="0000001010111000";
        when 3195 => y_in <= "10001100"; x_in <= "11111011"; z_correct<="0000001001000100";
        when 3196 => y_in <= "10001100"; x_in <= "11111100"; z_correct<="0000000111010000";
        when 3197 => y_in <= "10001100"; x_in <= "11111101"; z_correct<="0000000101011100";
        when 3198 => y_in <= "10001100"; x_in <= "11111110"; z_correct<="0000000011101000";
        when 3199 => y_in <= "10001100"; x_in <= "11111111"; z_correct<="0000000001110100";
        when 3200 => y_in <= "10001100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 3201 => y_in <= "10001100"; x_in <= "00000001"; z_correct<="1111111110001100";
        when 3202 => y_in <= "10001100"; x_in <= "00000010"; z_correct<="1111111100011000";
        when 3203 => y_in <= "10001100"; x_in <= "00000011"; z_correct<="1111111010100100";
        when 3204 => y_in <= "10001100"; x_in <= "00000100"; z_correct<="1111111000110000";
        when 3205 => y_in <= "10001100"; x_in <= "00000101"; z_correct<="1111110110111100";
        when 3206 => y_in <= "10001100"; x_in <= "00000110"; z_correct<="1111110101001000";
        when 3207 => y_in <= "10001100"; x_in <= "00000111"; z_correct<="1111110011010100";
        when 3208 => y_in <= "10001100"; x_in <= "00001000"; z_correct<="1111110001100000";
        when 3209 => y_in <= "10001100"; x_in <= "00001001"; z_correct<="1111101111101100";
        when 3210 => y_in <= "10001100"; x_in <= "00001010"; z_correct<="1111101101111000";
        when 3211 => y_in <= "10001100"; x_in <= "00001011"; z_correct<="1111101100000100";
        when 3212 => y_in <= "10001100"; x_in <= "00001100"; z_correct<="1111101010010000";
        when 3213 => y_in <= "10001100"; x_in <= "00001101"; z_correct<="1111101000011100";
        when 3214 => y_in <= "10001100"; x_in <= "00001110"; z_correct<="1111100110101000";
        when 3215 => y_in <= "10001100"; x_in <= "00001111"; z_correct<="1111100100110100";
        when 3216 => y_in <= "10001100"; x_in <= "00010000"; z_correct<="1111100011000000";
        when 3217 => y_in <= "10001100"; x_in <= "00010001"; z_correct<="1111100001001100";
        when 3218 => y_in <= "10001100"; x_in <= "00010010"; z_correct<="1111011111011000";
        when 3219 => y_in <= "10001100"; x_in <= "00010011"; z_correct<="1111011101100100";
        when 3220 => y_in <= "10001100"; x_in <= "00010100"; z_correct<="1111011011110000";
        when 3221 => y_in <= "10001100"; x_in <= "00010101"; z_correct<="1111011001111100";
        when 3222 => y_in <= "10001100"; x_in <= "00010110"; z_correct<="1111011000001000";
        when 3223 => y_in <= "10001100"; x_in <= "00010111"; z_correct<="1111010110010100";
        when 3224 => y_in <= "10001100"; x_in <= "00011000"; z_correct<="1111010100100000";
        when 3225 => y_in <= "10001100"; x_in <= "00011001"; z_correct<="1111010010101100";
        when 3226 => y_in <= "10001100"; x_in <= "00011010"; z_correct<="1111010000111000";
        when 3227 => y_in <= "10001100"; x_in <= "00011011"; z_correct<="1111001111000100";
        when 3228 => y_in <= "10001100"; x_in <= "00011100"; z_correct<="1111001101010000";
        when 3229 => y_in <= "10001100"; x_in <= "00011101"; z_correct<="1111001011011100";
        when 3230 => y_in <= "10001100"; x_in <= "00011110"; z_correct<="1111001001101000";
        when 3231 => y_in <= "10001100"; x_in <= "00011111"; z_correct<="1111000111110100";
        when 3232 => y_in <= "10001100"; x_in <= "00100000"; z_correct<="1111000110000000";
        when 3233 => y_in <= "10001100"; x_in <= "00100001"; z_correct<="1111000100001100";
        when 3234 => y_in <= "10001100"; x_in <= "00100010"; z_correct<="1111000010011000";
        when 3235 => y_in <= "10001100"; x_in <= "00100011"; z_correct<="1111000000100100";
        when 3236 => y_in <= "10001100"; x_in <= "00100100"; z_correct<="1110111110110000";
        when 3237 => y_in <= "10001100"; x_in <= "00100101"; z_correct<="1110111100111100";
        when 3238 => y_in <= "10001100"; x_in <= "00100110"; z_correct<="1110111011001000";
        when 3239 => y_in <= "10001100"; x_in <= "00100111"; z_correct<="1110111001010100";
        when 3240 => y_in <= "10001100"; x_in <= "00101000"; z_correct<="1110110111100000";
        when 3241 => y_in <= "10001100"; x_in <= "00101001"; z_correct<="1110110101101100";
        when 3242 => y_in <= "10001100"; x_in <= "00101010"; z_correct<="1110110011111000";
        when 3243 => y_in <= "10001100"; x_in <= "00101011"; z_correct<="1110110010000100";
        when 3244 => y_in <= "10001100"; x_in <= "00101100"; z_correct<="1110110000010000";
        when 3245 => y_in <= "10001100"; x_in <= "00101101"; z_correct<="1110101110011100";
        when 3246 => y_in <= "10001100"; x_in <= "00101110"; z_correct<="1110101100101000";
        when 3247 => y_in <= "10001100"; x_in <= "00101111"; z_correct<="1110101010110100";
        when 3248 => y_in <= "10001100"; x_in <= "00110000"; z_correct<="1110101001000000";
        when 3249 => y_in <= "10001100"; x_in <= "00110001"; z_correct<="1110100111001100";
        when 3250 => y_in <= "10001100"; x_in <= "00110010"; z_correct<="1110100101011000";
        when 3251 => y_in <= "10001100"; x_in <= "00110011"; z_correct<="1110100011100100";
        when 3252 => y_in <= "10001100"; x_in <= "00110100"; z_correct<="1110100001110000";
        when 3253 => y_in <= "10001100"; x_in <= "00110101"; z_correct<="1110011111111100";
        when 3254 => y_in <= "10001100"; x_in <= "00110110"; z_correct<="1110011110001000";
        when 3255 => y_in <= "10001100"; x_in <= "00110111"; z_correct<="1110011100010100";
        when 3256 => y_in <= "10001100"; x_in <= "00111000"; z_correct<="1110011010100000";
        when 3257 => y_in <= "10001100"; x_in <= "00111001"; z_correct<="1110011000101100";
        when 3258 => y_in <= "10001100"; x_in <= "00111010"; z_correct<="1110010110111000";
        when 3259 => y_in <= "10001100"; x_in <= "00111011"; z_correct<="1110010101000100";
        when 3260 => y_in <= "10001100"; x_in <= "00111100"; z_correct<="1110010011010000";
        when 3261 => y_in <= "10001100"; x_in <= "00111101"; z_correct<="1110010001011100";
        when 3262 => y_in <= "10001100"; x_in <= "00111110"; z_correct<="1110001111101000";
        when 3263 => y_in <= "10001100"; x_in <= "00111111"; z_correct<="1110001101110100";
        when 3264 => y_in <= "10001100"; x_in <= "01000000"; z_correct<="1110001100000000";
        when 3265 => y_in <= "10001100"; x_in <= "01000001"; z_correct<="1110001010001100";
        when 3266 => y_in <= "10001100"; x_in <= "01000010"; z_correct<="1110001000011000";
        when 3267 => y_in <= "10001100"; x_in <= "01000011"; z_correct<="1110000110100100";
        when 3268 => y_in <= "10001100"; x_in <= "01000100"; z_correct<="1110000100110000";
        when 3269 => y_in <= "10001100"; x_in <= "01000101"; z_correct<="1110000010111100";
        when 3270 => y_in <= "10001100"; x_in <= "01000110"; z_correct<="1110000001001000";
        when 3271 => y_in <= "10001100"; x_in <= "01000111"; z_correct<="1101111111010100";
        when 3272 => y_in <= "10001100"; x_in <= "01001000"; z_correct<="1101111101100000";
        when 3273 => y_in <= "10001100"; x_in <= "01001001"; z_correct<="1101111011101100";
        when 3274 => y_in <= "10001100"; x_in <= "01001010"; z_correct<="1101111001111000";
        when 3275 => y_in <= "10001100"; x_in <= "01001011"; z_correct<="1101111000000100";
        when 3276 => y_in <= "10001100"; x_in <= "01001100"; z_correct<="1101110110010000";
        when 3277 => y_in <= "10001100"; x_in <= "01001101"; z_correct<="1101110100011100";
        when 3278 => y_in <= "10001100"; x_in <= "01001110"; z_correct<="1101110010101000";
        when 3279 => y_in <= "10001100"; x_in <= "01001111"; z_correct<="1101110000110100";
        when 3280 => y_in <= "10001100"; x_in <= "01010000"; z_correct<="1101101111000000";
        when 3281 => y_in <= "10001100"; x_in <= "01010001"; z_correct<="1101101101001100";
        when 3282 => y_in <= "10001100"; x_in <= "01010010"; z_correct<="1101101011011000";
        when 3283 => y_in <= "10001100"; x_in <= "01010011"; z_correct<="1101101001100100";
        when 3284 => y_in <= "10001100"; x_in <= "01010100"; z_correct<="1101100111110000";
        when 3285 => y_in <= "10001100"; x_in <= "01010101"; z_correct<="1101100101111100";
        when 3286 => y_in <= "10001100"; x_in <= "01010110"; z_correct<="1101100100001000";
        when 3287 => y_in <= "10001100"; x_in <= "01010111"; z_correct<="1101100010010100";
        when 3288 => y_in <= "10001100"; x_in <= "01011000"; z_correct<="1101100000100000";
        when 3289 => y_in <= "10001100"; x_in <= "01011001"; z_correct<="1101011110101100";
        when 3290 => y_in <= "10001100"; x_in <= "01011010"; z_correct<="1101011100111000";
        when 3291 => y_in <= "10001100"; x_in <= "01011011"; z_correct<="1101011011000100";
        when 3292 => y_in <= "10001100"; x_in <= "01011100"; z_correct<="1101011001010000";
        when 3293 => y_in <= "10001100"; x_in <= "01011101"; z_correct<="1101010111011100";
        when 3294 => y_in <= "10001100"; x_in <= "01011110"; z_correct<="1101010101101000";
        when 3295 => y_in <= "10001100"; x_in <= "01011111"; z_correct<="1101010011110100";
        when 3296 => y_in <= "10001100"; x_in <= "01100000"; z_correct<="1101010010000000";
        when 3297 => y_in <= "10001100"; x_in <= "01100001"; z_correct<="1101010000001100";
        when 3298 => y_in <= "10001100"; x_in <= "01100010"; z_correct<="1101001110011000";
        when 3299 => y_in <= "10001100"; x_in <= "01100011"; z_correct<="1101001100100100";
        when 3300 => y_in <= "10001100"; x_in <= "01100100"; z_correct<="1101001010110000";
        when 3301 => y_in <= "10001100"; x_in <= "01100101"; z_correct<="1101001000111100";
        when 3302 => y_in <= "10001100"; x_in <= "01100110"; z_correct<="1101000111001000";
        when 3303 => y_in <= "10001100"; x_in <= "01100111"; z_correct<="1101000101010100";
        when 3304 => y_in <= "10001100"; x_in <= "01101000"; z_correct<="1101000011100000";
        when 3305 => y_in <= "10001100"; x_in <= "01101001"; z_correct<="1101000001101100";
        when 3306 => y_in <= "10001100"; x_in <= "01101010"; z_correct<="1100111111111000";
        when 3307 => y_in <= "10001100"; x_in <= "01101011"; z_correct<="1100111110000100";
        when 3308 => y_in <= "10001100"; x_in <= "01101100"; z_correct<="1100111100010000";
        when 3309 => y_in <= "10001100"; x_in <= "01101101"; z_correct<="1100111010011100";
        when 3310 => y_in <= "10001100"; x_in <= "01101110"; z_correct<="1100111000101000";
        when 3311 => y_in <= "10001100"; x_in <= "01101111"; z_correct<="1100110110110100";
        when 3312 => y_in <= "10001100"; x_in <= "01110000"; z_correct<="1100110101000000";
        when 3313 => y_in <= "10001100"; x_in <= "01110001"; z_correct<="1100110011001100";
        when 3314 => y_in <= "10001100"; x_in <= "01110010"; z_correct<="1100110001011000";
        when 3315 => y_in <= "10001100"; x_in <= "01110011"; z_correct<="1100101111100100";
        when 3316 => y_in <= "10001100"; x_in <= "01110100"; z_correct<="1100101101110000";
        when 3317 => y_in <= "10001100"; x_in <= "01110101"; z_correct<="1100101011111100";
        when 3318 => y_in <= "10001100"; x_in <= "01110110"; z_correct<="1100101010001000";
        when 3319 => y_in <= "10001100"; x_in <= "01110111"; z_correct<="1100101000010100";
        when 3320 => y_in <= "10001100"; x_in <= "01111000"; z_correct<="1100100110100000";
        when 3321 => y_in <= "10001100"; x_in <= "01111001"; z_correct<="1100100100101100";
        when 3322 => y_in <= "10001100"; x_in <= "01111010"; z_correct<="1100100010111000";
        when 3323 => y_in <= "10001100"; x_in <= "01111011"; z_correct<="1100100001000100";
        when 3324 => y_in <= "10001100"; x_in <= "01111100"; z_correct<="1100011111010000";
        when 3325 => y_in <= "10001100"; x_in <= "01111101"; z_correct<="1100011101011100";
        when 3326 => y_in <= "10001100"; x_in <= "01111110"; z_correct<="1100011011101000";
        when 3327 => y_in <= "10001100"; x_in <= "01111111"; z_correct<="1100011001110100";
        when 3328 => y_in <= "10001101"; x_in <= "10000000"; z_correct<="0011100110000000";
        when 3329 => y_in <= "10001101"; x_in <= "10000001"; z_correct<="0011100100001101";
        when 3330 => y_in <= "10001101"; x_in <= "10000010"; z_correct<="0011100010011010";
        when 3331 => y_in <= "10001101"; x_in <= "10000011"; z_correct<="0011100000100111";
        when 3332 => y_in <= "10001101"; x_in <= "10000100"; z_correct<="0011011110110100";
        when 3333 => y_in <= "10001101"; x_in <= "10000101"; z_correct<="0011011101000001";
        when 3334 => y_in <= "10001101"; x_in <= "10000110"; z_correct<="0011011011001110";
        when 3335 => y_in <= "10001101"; x_in <= "10000111"; z_correct<="0011011001011011";
        when 3336 => y_in <= "10001101"; x_in <= "10001000"; z_correct<="0011010111101000";
        when 3337 => y_in <= "10001101"; x_in <= "10001001"; z_correct<="0011010101110101";
        when 3338 => y_in <= "10001101"; x_in <= "10001010"; z_correct<="0011010100000010";
        when 3339 => y_in <= "10001101"; x_in <= "10001011"; z_correct<="0011010010001111";
        when 3340 => y_in <= "10001101"; x_in <= "10001100"; z_correct<="0011010000011100";
        when 3341 => y_in <= "10001101"; x_in <= "10001101"; z_correct<="0011001110101001";
        when 3342 => y_in <= "10001101"; x_in <= "10001110"; z_correct<="0011001100110110";
        when 3343 => y_in <= "10001101"; x_in <= "10001111"; z_correct<="0011001011000011";
        when 3344 => y_in <= "10001101"; x_in <= "10010000"; z_correct<="0011001001010000";
        when 3345 => y_in <= "10001101"; x_in <= "10010001"; z_correct<="0011000111011101";
        when 3346 => y_in <= "10001101"; x_in <= "10010010"; z_correct<="0011000101101010";
        when 3347 => y_in <= "10001101"; x_in <= "10010011"; z_correct<="0011000011110111";
        when 3348 => y_in <= "10001101"; x_in <= "10010100"; z_correct<="0011000010000100";
        when 3349 => y_in <= "10001101"; x_in <= "10010101"; z_correct<="0011000000010001";
        when 3350 => y_in <= "10001101"; x_in <= "10010110"; z_correct<="0010111110011110";
        when 3351 => y_in <= "10001101"; x_in <= "10010111"; z_correct<="0010111100101011";
        when 3352 => y_in <= "10001101"; x_in <= "10011000"; z_correct<="0010111010111000";
        when 3353 => y_in <= "10001101"; x_in <= "10011001"; z_correct<="0010111001000101";
        when 3354 => y_in <= "10001101"; x_in <= "10011010"; z_correct<="0010110111010010";
        when 3355 => y_in <= "10001101"; x_in <= "10011011"; z_correct<="0010110101011111";
        when 3356 => y_in <= "10001101"; x_in <= "10011100"; z_correct<="0010110011101100";
        when 3357 => y_in <= "10001101"; x_in <= "10011101"; z_correct<="0010110001111001";
        when 3358 => y_in <= "10001101"; x_in <= "10011110"; z_correct<="0010110000000110";
        when 3359 => y_in <= "10001101"; x_in <= "10011111"; z_correct<="0010101110010011";
        when 3360 => y_in <= "10001101"; x_in <= "10100000"; z_correct<="0010101100100000";
        when 3361 => y_in <= "10001101"; x_in <= "10100001"; z_correct<="0010101010101101";
        when 3362 => y_in <= "10001101"; x_in <= "10100010"; z_correct<="0010101000111010";
        when 3363 => y_in <= "10001101"; x_in <= "10100011"; z_correct<="0010100111000111";
        when 3364 => y_in <= "10001101"; x_in <= "10100100"; z_correct<="0010100101010100";
        when 3365 => y_in <= "10001101"; x_in <= "10100101"; z_correct<="0010100011100001";
        when 3366 => y_in <= "10001101"; x_in <= "10100110"; z_correct<="0010100001101110";
        when 3367 => y_in <= "10001101"; x_in <= "10100111"; z_correct<="0010011111111011";
        when 3368 => y_in <= "10001101"; x_in <= "10101000"; z_correct<="0010011110001000";
        when 3369 => y_in <= "10001101"; x_in <= "10101001"; z_correct<="0010011100010101";
        when 3370 => y_in <= "10001101"; x_in <= "10101010"; z_correct<="0010011010100010";
        when 3371 => y_in <= "10001101"; x_in <= "10101011"; z_correct<="0010011000101111";
        when 3372 => y_in <= "10001101"; x_in <= "10101100"; z_correct<="0010010110111100";
        when 3373 => y_in <= "10001101"; x_in <= "10101101"; z_correct<="0010010101001001";
        when 3374 => y_in <= "10001101"; x_in <= "10101110"; z_correct<="0010010011010110";
        when 3375 => y_in <= "10001101"; x_in <= "10101111"; z_correct<="0010010001100011";
        when 3376 => y_in <= "10001101"; x_in <= "10110000"; z_correct<="0010001111110000";
        when 3377 => y_in <= "10001101"; x_in <= "10110001"; z_correct<="0010001101111101";
        when 3378 => y_in <= "10001101"; x_in <= "10110010"; z_correct<="0010001100001010";
        when 3379 => y_in <= "10001101"; x_in <= "10110011"; z_correct<="0010001010010111";
        when 3380 => y_in <= "10001101"; x_in <= "10110100"; z_correct<="0010001000100100";
        when 3381 => y_in <= "10001101"; x_in <= "10110101"; z_correct<="0010000110110001";
        when 3382 => y_in <= "10001101"; x_in <= "10110110"; z_correct<="0010000100111110";
        when 3383 => y_in <= "10001101"; x_in <= "10110111"; z_correct<="0010000011001011";
        when 3384 => y_in <= "10001101"; x_in <= "10111000"; z_correct<="0010000001011000";
        when 3385 => y_in <= "10001101"; x_in <= "10111001"; z_correct<="0001111111100101";
        when 3386 => y_in <= "10001101"; x_in <= "10111010"; z_correct<="0001111101110010";
        when 3387 => y_in <= "10001101"; x_in <= "10111011"; z_correct<="0001111011111111";
        when 3388 => y_in <= "10001101"; x_in <= "10111100"; z_correct<="0001111010001100";
        when 3389 => y_in <= "10001101"; x_in <= "10111101"; z_correct<="0001111000011001";
        when 3390 => y_in <= "10001101"; x_in <= "10111110"; z_correct<="0001110110100110";
        when 3391 => y_in <= "10001101"; x_in <= "10111111"; z_correct<="0001110100110011";
        when 3392 => y_in <= "10001101"; x_in <= "11000000"; z_correct<="0001110011000000";
        when 3393 => y_in <= "10001101"; x_in <= "11000001"; z_correct<="0001110001001101";
        when 3394 => y_in <= "10001101"; x_in <= "11000010"; z_correct<="0001101111011010";
        when 3395 => y_in <= "10001101"; x_in <= "11000011"; z_correct<="0001101101100111";
        when 3396 => y_in <= "10001101"; x_in <= "11000100"; z_correct<="0001101011110100";
        when 3397 => y_in <= "10001101"; x_in <= "11000101"; z_correct<="0001101010000001";
        when 3398 => y_in <= "10001101"; x_in <= "11000110"; z_correct<="0001101000001110";
        when 3399 => y_in <= "10001101"; x_in <= "11000111"; z_correct<="0001100110011011";
        when 3400 => y_in <= "10001101"; x_in <= "11001000"; z_correct<="0001100100101000";
        when 3401 => y_in <= "10001101"; x_in <= "11001001"; z_correct<="0001100010110101";
        when 3402 => y_in <= "10001101"; x_in <= "11001010"; z_correct<="0001100001000010";
        when 3403 => y_in <= "10001101"; x_in <= "11001011"; z_correct<="0001011111001111";
        when 3404 => y_in <= "10001101"; x_in <= "11001100"; z_correct<="0001011101011100";
        when 3405 => y_in <= "10001101"; x_in <= "11001101"; z_correct<="0001011011101001";
        when 3406 => y_in <= "10001101"; x_in <= "11001110"; z_correct<="0001011001110110";
        when 3407 => y_in <= "10001101"; x_in <= "11001111"; z_correct<="0001011000000011";
        when 3408 => y_in <= "10001101"; x_in <= "11010000"; z_correct<="0001010110010000";
        when 3409 => y_in <= "10001101"; x_in <= "11010001"; z_correct<="0001010100011101";
        when 3410 => y_in <= "10001101"; x_in <= "11010010"; z_correct<="0001010010101010";
        when 3411 => y_in <= "10001101"; x_in <= "11010011"; z_correct<="0001010000110111";
        when 3412 => y_in <= "10001101"; x_in <= "11010100"; z_correct<="0001001111000100";
        when 3413 => y_in <= "10001101"; x_in <= "11010101"; z_correct<="0001001101010001";
        when 3414 => y_in <= "10001101"; x_in <= "11010110"; z_correct<="0001001011011110";
        when 3415 => y_in <= "10001101"; x_in <= "11010111"; z_correct<="0001001001101011";
        when 3416 => y_in <= "10001101"; x_in <= "11011000"; z_correct<="0001000111111000";
        when 3417 => y_in <= "10001101"; x_in <= "11011001"; z_correct<="0001000110000101";
        when 3418 => y_in <= "10001101"; x_in <= "11011010"; z_correct<="0001000100010010";
        when 3419 => y_in <= "10001101"; x_in <= "11011011"; z_correct<="0001000010011111";
        when 3420 => y_in <= "10001101"; x_in <= "11011100"; z_correct<="0001000000101100";
        when 3421 => y_in <= "10001101"; x_in <= "11011101"; z_correct<="0000111110111001";
        when 3422 => y_in <= "10001101"; x_in <= "11011110"; z_correct<="0000111101000110";
        when 3423 => y_in <= "10001101"; x_in <= "11011111"; z_correct<="0000111011010011";
        when 3424 => y_in <= "10001101"; x_in <= "11100000"; z_correct<="0000111001100000";
        when 3425 => y_in <= "10001101"; x_in <= "11100001"; z_correct<="0000110111101101";
        when 3426 => y_in <= "10001101"; x_in <= "11100010"; z_correct<="0000110101111010";
        when 3427 => y_in <= "10001101"; x_in <= "11100011"; z_correct<="0000110100000111";
        when 3428 => y_in <= "10001101"; x_in <= "11100100"; z_correct<="0000110010010100";
        when 3429 => y_in <= "10001101"; x_in <= "11100101"; z_correct<="0000110000100001";
        when 3430 => y_in <= "10001101"; x_in <= "11100110"; z_correct<="0000101110101110";
        when 3431 => y_in <= "10001101"; x_in <= "11100111"; z_correct<="0000101100111011";
        when 3432 => y_in <= "10001101"; x_in <= "11101000"; z_correct<="0000101011001000";
        when 3433 => y_in <= "10001101"; x_in <= "11101001"; z_correct<="0000101001010101";
        when 3434 => y_in <= "10001101"; x_in <= "11101010"; z_correct<="0000100111100010";
        when 3435 => y_in <= "10001101"; x_in <= "11101011"; z_correct<="0000100101101111";
        when 3436 => y_in <= "10001101"; x_in <= "11101100"; z_correct<="0000100011111100";
        when 3437 => y_in <= "10001101"; x_in <= "11101101"; z_correct<="0000100010001001";
        when 3438 => y_in <= "10001101"; x_in <= "11101110"; z_correct<="0000100000010110";
        when 3439 => y_in <= "10001101"; x_in <= "11101111"; z_correct<="0000011110100011";
        when 3440 => y_in <= "10001101"; x_in <= "11110000"; z_correct<="0000011100110000";
        when 3441 => y_in <= "10001101"; x_in <= "11110001"; z_correct<="0000011010111101";
        when 3442 => y_in <= "10001101"; x_in <= "11110010"; z_correct<="0000011001001010";
        when 3443 => y_in <= "10001101"; x_in <= "11110011"; z_correct<="0000010111010111";
        when 3444 => y_in <= "10001101"; x_in <= "11110100"; z_correct<="0000010101100100";
        when 3445 => y_in <= "10001101"; x_in <= "11110101"; z_correct<="0000010011110001";
        when 3446 => y_in <= "10001101"; x_in <= "11110110"; z_correct<="0000010001111110";
        when 3447 => y_in <= "10001101"; x_in <= "11110111"; z_correct<="0000010000001011";
        when 3448 => y_in <= "10001101"; x_in <= "11111000"; z_correct<="0000001110011000";
        when 3449 => y_in <= "10001101"; x_in <= "11111001"; z_correct<="0000001100100101";
        when 3450 => y_in <= "10001101"; x_in <= "11111010"; z_correct<="0000001010110010";
        when 3451 => y_in <= "10001101"; x_in <= "11111011"; z_correct<="0000001000111111";
        when 3452 => y_in <= "10001101"; x_in <= "11111100"; z_correct<="0000000111001100";
        when 3453 => y_in <= "10001101"; x_in <= "11111101"; z_correct<="0000000101011001";
        when 3454 => y_in <= "10001101"; x_in <= "11111110"; z_correct<="0000000011100110";
        when 3455 => y_in <= "10001101"; x_in <= "11111111"; z_correct<="0000000001110011";
        when 3456 => y_in <= "10001101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 3457 => y_in <= "10001101"; x_in <= "00000001"; z_correct<="1111111110001101";
        when 3458 => y_in <= "10001101"; x_in <= "00000010"; z_correct<="1111111100011010";
        when 3459 => y_in <= "10001101"; x_in <= "00000011"; z_correct<="1111111010100111";
        when 3460 => y_in <= "10001101"; x_in <= "00000100"; z_correct<="1111111000110100";
        when 3461 => y_in <= "10001101"; x_in <= "00000101"; z_correct<="1111110111000001";
        when 3462 => y_in <= "10001101"; x_in <= "00000110"; z_correct<="1111110101001110";
        when 3463 => y_in <= "10001101"; x_in <= "00000111"; z_correct<="1111110011011011";
        when 3464 => y_in <= "10001101"; x_in <= "00001000"; z_correct<="1111110001101000";
        when 3465 => y_in <= "10001101"; x_in <= "00001001"; z_correct<="1111101111110101";
        when 3466 => y_in <= "10001101"; x_in <= "00001010"; z_correct<="1111101110000010";
        when 3467 => y_in <= "10001101"; x_in <= "00001011"; z_correct<="1111101100001111";
        when 3468 => y_in <= "10001101"; x_in <= "00001100"; z_correct<="1111101010011100";
        when 3469 => y_in <= "10001101"; x_in <= "00001101"; z_correct<="1111101000101001";
        when 3470 => y_in <= "10001101"; x_in <= "00001110"; z_correct<="1111100110110110";
        when 3471 => y_in <= "10001101"; x_in <= "00001111"; z_correct<="1111100101000011";
        when 3472 => y_in <= "10001101"; x_in <= "00010000"; z_correct<="1111100011010000";
        when 3473 => y_in <= "10001101"; x_in <= "00010001"; z_correct<="1111100001011101";
        when 3474 => y_in <= "10001101"; x_in <= "00010010"; z_correct<="1111011111101010";
        when 3475 => y_in <= "10001101"; x_in <= "00010011"; z_correct<="1111011101110111";
        when 3476 => y_in <= "10001101"; x_in <= "00010100"; z_correct<="1111011100000100";
        when 3477 => y_in <= "10001101"; x_in <= "00010101"; z_correct<="1111011010010001";
        when 3478 => y_in <= "10001101"; x_in <= "00010110"; z_correct<="1111011000011110";
        when 3479 => y_in <= "10001101"; x_in <= "00010111"; z_correct<="1111010110101011";
        when 3480 => y_in <= "10001101"; x_in <= "00011000"; z_correct<="1111010100111000";
        when 3481 => y_in <= "10001101"; x_in <= "00011001"; z_correct<="1111010011000101";
        when 3482 => y_in <= "10001101"; x_in <= "00011010"; z_correct<="1111010001010010";
        when 3483 => y_in <= "10001101"; x_in <= "00011011"; z_correct<="1111001111011111";
        when 3484 => y_in <= "10001101"; x_in <= "00011100"; z_correct<="1111001101101100";
        when 3485 => y_in <= "10001101"; x_in <= "00011101"; z_correct<="1111001011111001";
        when 3486 => y_in <= "10001101"; x_in <= "00011110"; z_correct<="1111001010000110";
        when 3487 => y_in <= "10001101"; x_in <= "00011111"; z_correct<="1111001000010011";
        when 3488 => y_in <= "10001101"; x_in <= "00100000"; z_correct<="1111000110100000";
        when 3489 => y_in <= "10001101"; x_in <= "00100001"; z_correct<="1111000100101101";
        when 3490 => y_in <= "10001101"; x_in <= "00100010"; z_correct<="1111000010111010";
        when 3491 => y_in <= "10001101"; x_in <= "00100011"; z_correct<="1111000001000111";
        when 3492 => y_in <= "10001101"; x_in <= "00100100"; z_correct<="1110111111010100";
        when 3493 => y_in <= "10001101"; x_in <= "00100101"; z_correct<="1110111101100001";
        when 3494 => y_in <= "10001101"; x_in <= "00100110"; z_correct<="1110111011101110";
        when 3495 => y_in <= "10001101"; x_in <= "00100111"; z_correct<="1110111001111011";
        when 3496 => y_in <= "10001101"; x_in <= "00101000"; z_correct<="1110111000001000";
        when 3497 => y_in <= "10001101"; x_in <= "00101001"; z_correct<="1110110110010101";
        when 3498 => y_in <= "10001101"; x_in <= "00101010"; z_correct<="1110110100100010";
        when 3499 => y_in <= "10001101"; x_in <= "00101011"; z_correct<="1110110010101111";
        when 3500 => y_in <= "10001101"; x_in <= "00101100"; z_correct<="1110110000111100";
        when 3501 => y_in <= "10001101"; x_in <= "00101101"; z_correct<="1110101111001001";
        when 3502 => y_in <= "10001101"; x_in <= "00101110"; z_correct<="1110101101010110";
        when 3503 => y_in <= "10001101"; x_in <= "00101111"; z_correct<="1110101011100011";
        when 3504 => y_in <= "10001101"; x_in <= "00110000"; z_correct<="1110101001110000";
        when 3505 => y_in <= "10001101"; x_in <= "00110001"; z_correct<="1110100111111101";
        when 3506 => y_in <= "10001101"; x_in <= "00110010"; z_correct<="1110100110001010";
        when 3507 => y_in <= "10001101"; x_in <= "00110011"; z_correct<="1110100100010111";
        when 3508 => y_in <= "10001101"; x_in <= "00110100"; z_correct<="1110100010100100";
        when 3509 => y_in <= "10001101"; x_in <= "00110101"; z_correct<="1110100000110001";
        when 3510 => y_in <= "10001101"; x_in <= "00110110"; z_correct<="1110011110111110";
        when 3511 => y_in <= "10001101"; x_in <= "00110111"; z_correct<="1110011101001011";
        when 3512 => y_in <= "10001101"; x_in <= "00111000"; z_correct<="1110011011011000";
        when 3513 => y_in <= "10001101"; x_in <= "00111001"; z_correct<="1110011001100101";
        when 3514 => y_in <= "10001101"; x_in <= "00111010"; z_correct<="1110010111110010";
        when 3515 => y_in <= "10001101"; x_in <= "00111011"; z_correct<="1110010101111111";
        when 3516 => y_in <= "10001101"; x_in <= "00111100"; z_correct<="1110010100001100";
        when 3517 => y_in <= "10001101"; x_in <= "00111101"; z_correct<="1110010010011001";
        when 3518 => y_in <= "10001101"; x_in <= "00111110"; z_correct<="1110010000100110";
        when 3519 => y_in <= "10001101"; x_in <= "00111111"; z_correct<="1110001110110011";
        when 3520 => y_in <= "10001101"; x_in <= "01000000"; z_correct<="1110001101000000";
        when 3521 => y_in <= "10001101"; x_in <= "01000001"; z_correct<="1110001011001101";
        when 3522 => y_in <= "10001101"; x_in <= "01000010"; z_correct<="1110001001011010";
        when 3523 => y_in <= "10001101"; x_in <= "01000011"; z_correct<="1110000111100111";
        when 3524 => y_in <= "10001101"; x_in <= "01000100"; z_correct<="1110000101110100";
        when 3525 => y_in <= "10001101"; x_in <= "01000101"; z_correct<="1110000100000001";
        when 3526 => y_in <= "10001101"; x_in <= "01000110"; z_correct<="1110000010001110";
        when 3527 => y_in <= "10001101"; x_in <= "01000111"; z_correct<="1110000000011011";
        when 3528 => y_in <= "10001101"; x_in <= "01001000"; z_correct<="1101111110101000";
        when 3529 => y_in <= "10001101"; x_in <= "01001001"; z_correct<="1101111100110101";
        when 3530 => y_in <= "10001101"; x_in <= "01001010"; z_correct<="1101111011000010";
        when 3531 => y_in <= "10001101"; x_in <= "01001011"; z_correct<="1101111001001111";
        when 3532 => y_in <= "10001101"; x_in <= "01001100"; z_correct<="1101110111011100";
        when 3533 => y_in <= "10001101"; x_in <= "01001101"; z_correct<="1101110101101001";
        when 3534 => y_in <= "10001101"; x_in <= "01001110"; z_correct<="1101110011110110";
        when 3535 => y_in <= "10001101"; x_in <= "01001111"; z_correct<="1101110010000011";
        when 3536 => y_in <= "10001101"; x_in <= "01010000"; z_correct<="1101110000010000";
        when 3537 => y_in <= "10001101"; x_in <= "01010001"; z_correct<="1101101110011101";
        when 3538 => y_in <= "10001101"; x_in <= "01010010"; z_correct<="1101101100101010";
        when 3539 => y_in <= "10001101"; x_in <= "01010011"; z_correct<="1101101010110111";
        when 3540 => y_in <= "10001101"; x_in <= "01010100"; z_correct<="1101101001000100";
        when 3541 => y_in <= "10001101"; x_in <= "01010101"; z_correct<="1101100111010001";
        when 3542 => y_in <= "10001101"; x_in <= "01010110"; z_correct<="1101100101011110";
        when 3543 => y_in <= "10001101"; x_in <= "01010111"; z_correct<="1101100011101011";
        when 3544 => y_in <= "10001101"; x_in <= "01011000"; z_correct<="1101100001111000";
        when 3545 => y_in <= "10001101"; x_in <= "01011001"; z_correct<="1101100000000101";
        when 3546 => y_in <= "10001101"; x_in <= "01011010"; z_correct<="1101011110010010";
        when 3547 => y_in <= "10001101"; x_in <= "01011011"; z_correct<="1101011100011111";
        when 3548 => y_in <= "10001101"; x_in <= "01011100"; z_correct<="1101011010101100";
        when 3549 => y_in <= "10001101"; x_in <= "01011101"; z_correct<="1101011000111001";
        when 3550 => y_in <= "10001101"; x_in <= "01011110"; z_correct<="1101010111000110";
        when 3551 => y_in <= "10001101"; x_in <= "01011111"; z_correct<="1101010101010011";
        when 3552 => y_in <= "10001101"; x_in <= "01100000"; z_correct<="1101010011100000";
        when 3553 => y_in <= "10001101"; x_in <= "01100001"; z_correct<="1101010001101101";
        when 3554 => y_in <= "10001101"; x_in <= "01100010"; z_correct<="1101001111111010";
        when 3555 => y_in <= "10001101"; x_in <= "01100011"; z_correct<="1101001110000111";
        when 3556 => y_in <= "10001101"; x_in <= "01100100"; z_correct<="1101001100010100";
        when 3557 => y_in <= "10001101"; x_in <= "01100101"; z_correct<="1101001010100001";
        when 3558 => y_in <= "10001101"; x_in <= "01100110"; z_correct<="1101001000101110";
        when 3559 => y_in <= "10001101"; x_in <= "01100111"; z_correct<="1101000110111011";
        when 3560 => y_in <= "10001101"; x_in <= "01101000"; z_correct<="1101000101001000";
        when 3561 => y_in <= "10001101"; x_in <= "01101001"; z_correct<="1101000011010101";
        when 3562 => y_in <= "10001101"; x_in <= "01101010"; z_correct<="1101000001100010";
        when 3563 => y_in <= "10001101"; x_in <= "01101011"; z_correct<="1100111111101111";
        when 3564 => y_in <= "10001101"; x_in <= "01101100"; z_correct<="1100111101111100";
        when 3565 => y_in <= "10001101"; x_in <= "01101101"; z_correct<="1100111100001001";
        when 3566 => y_in <= "10001101"; x_in <= "01101110"; z_correct<="1100111010010110";
        when 3567 => y_in <= "10001101"; x_in <= "01101111"; z_correct<="1100111000100011";
        when 3568 => y_in <= "10001101"; x_in <= "01110000"; z_correct<="1100110110110000";
        when 3569 => y_in <= "10001101"; x_in <= "01110001"; z_correct<="1100110100111101";
        when 3570 => y_in <= "10001101"; x_in <= "01110010"; z_correct<="1100110011001010";
        when 3571 => y_in <= "10001101"; x_in <= "01110011"; z_correct<="1100110001010111";
        when 3572 => y_in <= "10001101"; x_in <= "01110100"; z_correct<="1100101111100100";
        when 3573 => y_in <= "10001101"; x_in <= "01110101"; z_correct<="1100101101110001";
        when 3574 => y_in <= "10001101"; x_in <= "01110110"; z_correct<="1100101011111110";
        when 3575 => y_in <= "10001101"; x_in <= "01110111"; z_correct<="1100101010001011";
        when 3576 => y_in <= "10001101"; x_in <= "01111000"; z_correct<="1100101000011000";
        when 3577 => y_in <= "10001101"; x_in <= "01111001"; z_correct<="1100100110100101";
        when 3578 => y_in <= "10001101"; x_in <= "01111010"; z_correct<="1100100100110010";
        when 3579 => y_in <= "10001101"; x_in <= "01111011"; z_correct<="1100100010111111";
        when 3580 => y_in <= "10001101"; x_in <= "01111100"; z_correct<="1100100001001100";
        when 3581 => y_in <= "10001101"; x_in <= "01111101"; z_correct<="1100011111011001";
        when 3582 => y_in <= "10001101"; x_in <= "01111110"; z_correct<="1100011101100110";
        when 3583 => y_in <= "10001101"; x_in <= "01111111"; z_correct<="1100011011110011";
        when 3584 => y_in <= "10001110"; x_in <= "10000000"; z_correct<="0011100100000000";
        when 3585 => y_in <= "10001110"; x_in <= "10000001"; z_correct<="0011100010001110";
        when 3586 => y_in <= "10001110"; x_in <= "10000010"; z_correct<="0011100000011100";
        when 3587 => y_in <= "10001110"; x_in <= "10000011"; z_correct<="0011011110101010";
        when 3588 => y_in <= "10001110"; x_in <= "10000100"; z_correct<="0011011100111000";
        when 3589 => y_in <= "10001110"; x_in <= "10000101"; z_correct<="0011011011000110";
        when 3590 => y_in <= "10001110"; x_in <= "10000110"; z_correct<="0011011001010100";
        when 3591 => y_in <= "10001110"; x_in <= "10000111"; z_correct<="0011010111100010";
        when 3592 => y_in <= "10001110"; x_in <= "10001000"; z_correct<="0011010101110000";
        when 3593 => y_in <= "10001110"; x_in <= "10001001"; z_correct<="0011010011111110";
        when 3594 => y_in <= "10001110"; x_in <= "10001010"; z_correct<="0011010010001100";
        when 3595 => y_in <= "10001110"; x_in <= "10001011"; z_correct<="0011010000011010";
        when 3596 => y_in <= "10001110"; x_in <= "10001100"; z_correct<="0011001110101000";
        when 3597 => y_in <= "10001110"; x_in <= "10001101"; z_correct<="0011001100110110";
        when 3598 => y_in <= "10001110"; x_in <= "10001110"; z_correct<="0011001011000100";
        when 3599 => y_in <= "10001110"; x_in <= "10001111"; z_correct<="0011001001010010";
        when 3600 => y_in <= "10001110"; x_in <= "10010000"; z_correct<="0011000111100000";
        when 3601 => y_in <= "10001110"; x_in <= "10010001"; z_correct<="0011000101101110";
        when 3602 => y_in <= "10001110"; x_in <= "10010010"; z_correct<="0011000011111100";
        when 3603 => y_in <= "10001110"; x_in <= "10010011"; z_correct<="0011000010001010";
        when 3604 => y_in <= "10001110"; x_in <= "10010100"; z_correct<="0011000000011000";
        when 3605 => y_in <= "10001110"; x_in <= "10010101"; z_correct<="0010111110100110";
        when 3606 => y_in <= "10001110"; x_in <= "10010110"; z_correct<="0010111100110100";
        when 3607 => y_in <= "10001110"; x_in <= "10010111"; z_correct<="0010111011000010";
        when 3608 => y_in <= "10001110"; x_in <= "10011000"; z_correct<="0010111001010000";
        when 3609 => y_in <= "10001110"; x_in <= "10011001"; z_correct<="0010110111011110";
        when 3610 => y_in <= "10001110"; x_in <= "10011010"; z_correct<="0010110101101100";
        when 3611 => y_in <= "10001110"; x_in <= "10011011"; z_correct<="0010110011111010";
        when 3612 => y_in <= "10001110"; x_in <= "10011100"; z_correct<="0010110010001000";
        when 3613 => y_in <= "10001110"; x_in <= "10011101"; z_correct<="0010110000010110";
        when 3614 => y_in <= "10001110"; x_in <= "10011110"; z_correct<="0010101110100100";
        when 3615 => y_in <= "10001110"; x_in <= "10011111"; z_correct<="0010101100110010";
        when 3616 => y_in <= "10001110"; x_in <= "10100000"; z_correct<="0010101011000000";
        when 3617 => y_in <= "10001110"; x_in <= "10100001"; z_correct<="0010101001001110";
        when 3618 => y_in <= "10001110"; x_in <= "10100010"; z_correct<="0010100111011100";
        when 3619 => y_in <= "10001110"; x_in <= "10100011"; z_correct<="0010100101101010";
        when 3620 => y_in <= "10001110"; x_in <= "10100100"; z_correct<="0010100011111000";
        when 3621 => y_in <= "10001110"; x_in <= "10100101"; z_correct<="0010100010000110";
        when 3622 => y_in <= "10001110"; x_in <= "10100110"; z_correct<="0010100000010100";
        when 3623 => y_in <= "10001110"; x_in <= "10100111"; z_correct<="0010011110100010";
        when 3624 => y_in <= "10001110"; x_in <= "10101000"; z_correct<="0010011100110000";
        when 3625 => y_in <= "10001110"; x_in <= "10101001"; z_correct<="0010011010111110";
        when 3626 => y_in <= "10001110"; x_in <= "10101010"; z_correct<="0010011001001100";
        when 3627 => y_in <= "10001110"; x_in <= "10101011"; z_correct<="0010010111011010";
        when 3628 => y_in <= "10001110"; x_in <= "10101100"; z_correct<="0010010101101000";
        when 3629 => y_in <= "10001110"; x_in <= "10101101"; z_correct<="0010010011110110";
        when 3630 => y_in <= "10001110"; x_in <= "10101110"; z_correct<="0010010010000100";
        when 3631 => y_in <= "10001110"; x_in <= "10101111"; z_correct<="0010010000010010";
        when 3632 => y_in <= "10001110"; x_in <= "10110000"; z_correct<="0010001110100000";
        when 3633 => y_in <= "10001110"; x_in <= "10110001"; z_correct<="0010001100101110";
        when 3634 => y_in <= "10001110"; x_in <= "10110010"; z_correct<="0010001010111100";
        when 3635 => y_in <= "10001110"; x_in <= "10110011"; z_correct<="0010001001001010";
        when 3636 => y_in <= "10001110"; x_in <= "10110100"; z_correct<="0010000111011000";
        when 3637 => y_in <= "10001110"; x_in <= "10110101"; z_correct<="0010000101100110";
        when 3638 => y_in <= "10001110"; x_in <= "10110110"; z_correct<="0010000011110100";
        when 3639 => y_in <= "10001110"; x_in <= "10110111"; z_correct<="0010000010000010";
        when 3640 => y_in <= "10001110"; x_in <= "10111000"; z_correct<="0010000000010000";
        when 3641 => y_in <= "10001110"; x_in <= "10111001"; z_correct<="0001111110011110";
        when 3642 => y_in <= "10001110"; x_in <= "10111010"; z_correct<="0001111100101100";
        when 3643 => y_in <= "10001110"; x_in <= "10111011"; z_correct<="0001111010111010";
        when 3644 => y_in <= "10001110"; x_in <= "10111100"; z_correct<="0001111001001000";
        when 3645 => y_in <= "10001110"; x_in <= "10111101"; z_correct<="0001110111010110";
        when 3646 => y_in <= "10001110"; x_in <= "10111110"; z_correct<="0001110101100100";
        when 3647 => y_in <= "10001110"; x_in <= "10111111"; z_correct<="0001110011110010";
        when 3648 => y_in <= "10001110"; x_in <= "11000000"; z_correct<="0001110010000000";
        when 3649 => y_in <= "10001110"; x_in <= "11000001"; z_correct<="0001110000001110";
        when 3650 => y_in <= "10001110"; x_in <= "11000010"; z_correct<="0001101110011100";
        when 3651 => y_in <= "10001110"; x_in <= "11000011"; z_correct<="0001101100101010";
        when 3652 => y_in <= "10001110"; x_in <= "11000100"; z_correct<="0001101010111000";
        when 3653 => y_in <= "10001110"; x_in <= "11000101"; z_correct<="0001101001000110";
        when 3654 => y_in <= "10001110"; x_in <= "11000110"; z_correct<="0001100111010100";
        when 3655 => y_in <= "10001110"; x_in <= "11000111"; z_correct<="0001100101100010";
        when 3656 => y_in <= "10001110"; x_in <= "11001000"; z_correct<="0001100011110000";
        when 3657 => y_in <= "10001110"; x_in <= "11001001"; z_correct<="0001100001111110";
        when 3658 => y_in <= "10001110"; x_in <= "11001010"; z_correct<="0001100000001100";
        when 3659 => y_in <= "10001110"; x_in <= "11001011"; z_correct<="0001011110011010";
        when 3660 => y_in <= "10001110"; x_in <= "11001100"; z_correct<="0001011100101000";
        when 3661 => y_in <= "10001110"; x_in <= "11001101"; z_correct<="0001011010110110";
        when 3662 => y_in <= "10001110"; x_in <= "11001110"; z_correct<="0001011001000100";
        when 3663 => y_in <= "10001110"; x_in <= "11001111"; z_correct<="0001010111010010";
        when 3664 => y_in <= "10001110"; x_in <= "11010000"; z_correct<="0001010101100000";
        when 3665 => y_in <= "10001110"; x_in <= "11010001"; z_correct<="0001010011101110";
        when 3666 => y_in <= "10001110"; x_in <= "11010010"; z_correct<="0001010001111100";
        when 3667 => y_in <= "10001110"; x_in <= "11010011"; z_correct<="0001010000001010";
        when 3668 => y_in <= "10001110"; x_in <= "11010100"; z_correct<="0001001110011000";
        when 3669 => y_in <= "10001110"; x_in <= "11010101"; z_correct<="0001001100100110";
        when 3670 => y_in <= "10001110"; x_in <= "11010110"; z_correct<="0001001010110100";
        when 3671 => y_in <= "10001110"; x_in <= "11010111"; z_correct<="0001001001000010";
        when 3672 => y_in <= "10001110"; x_in <= "11011000"; z_correct<="0001000111010000";
        when 3673 => y_in <= "10001110"; x_in <= "11011001"; z_correct<="0001000101011110";
        when 3674 => y_in <= "10001110"; x_in <= "11011010"; z_correct<="0001000011101100";
        when 3675 => y_in <= "10001110"; x_in <= "11011011"; z_correct<="0001000001111010";
        when 3676 => y_in <= "10001110"; x_in <= "11011100"; z_correct<="0001000000001000";
        when 3677 => y_in <= "10001110"; x_in <= "11011101"; z_correct<="0000111110010110";
        when 3678 => y_in <= "10001110"; x_in <= "11011110"; z_correct<="0000111100100100";
        when 3679 => y_in <= "10001110"; x_in <= "11011111"; z_correct<="0000111010110010";
        when 3680 => y_in <= "10001110"; x_in <= "11100000"; z_correct<="0000111001000000";
        when 3681 => y_in <= "10001110"; x_in <= "11100001"; z_correct<="0000110111001110";
        when 3682 => y_in <= "10001110"; x_in <= "11100010"; z_correct<="0000110101011100";
        when 3683 => y_in <= "10001110"; x_in <= "11100011"; z_correct<="0000110011101010";
        when 3684 => y_in <= "10001110"; x_in <= "11100100"; z_correct<="0000110001111000";
        when 3685 => y_in <= "10001110"; x_in <= "11100101"; z_correct<="0000110000000110";
        when 3686 => y_in <= "10001110"; x_in <= "11100110"; z_correct<="0000101110010100";
        when 3687 => y_in <= "10001110"; x_in <= "11100111"; z_correct<="0000101100100010";
        when 3688 => y_in <= "10001110"; x_in <= "11101000"; z_correct<="0000101010110000";
        when 3689 => y_in <= "10001110"; x_in <= "11101001"; z_correct<="0000101000111110";
        when 3690 => y_in <= "10001110"; x_in <= "11101010"; z_correct<="0000100111001100";
        when 3691 => y_in <= "10001110"; x_in <= "11101011"; z_correct<="0000100101011010";
        when 3692 => y_in <= "10001110"; x_in <= "11101100"; z_correct<="0000100011101000";
        when 3693 => y_in <= "10001110"; x_in <= "11101101"; z_correct<="0000100001110110";
        when 3694 => y_in <= "10001110"; x_in <= "11101110"; z_correct<="0000100000000100";
        when 3695 => y_in <= "10001110"; x_in <= "11101111"; z_correct<="0000011110010010";
        when 3696 => y_in <= "10001110"; x_in <= "11110000"; z_correct<="0000011100100000";
        when 3697 => y_in <= "10001110"; x_in <= "11110001"; z_correct<="0000011010101110";
        when 3698 => y_in <= "10001110"; x_in <= "11110010"; z_correct<="0000011000111100";
        when 3699 => y_in <= "10001110"; x_in <= "11110011"; z_correct<="0000010111001010";
        when 3700 => y_in <= "10001110"; x_in <= "11110100"; z_correct<="0000010101011000";
        when 3701 => y_in <= "10001110"; x_in <= "11110101"; z_correct<="0000010011100110";
        when 3702 => y_in <= "10001110"; x_in <= "11110110"; z_correct<="0000010001110100";
        when 3703 => y_in <= "10001110"; x_in <= "11110111"; z_correct<="0000010000000010";
        when 3704 => y_in <= "10001110"; x_in <= "11111000"; z_correct<="0000001110010000";
        when 3705 => y_in <= "10001110"; x_in <= "11111001"; z_correct<="0000001100011110";
        when 3706 => y_in <= "10001110"; x_in <= "11111010"; z_correct<="0000001010101100";
        when 3707 => y_in <= "10001110"; x_in <= "11111011"; z_correct<="0000001000111010";
        when 3708 => y_in <= "10001110"; x_in <= "11111100"; z_correct<="0000000111001000";
        when 3709 => y_in <= "10001110"; x_in <= "11111101"; z_correct<="0000000101010110";
        when 3710 => y_in <= "10001110"; x_in <= "11111110"; z_correct<="0000000011100100";
        when 3711 => y_in <= "10001110"; x_in <= "11111111"; z_correct<="0000000001110010";
        when 3712 => y_in <= "10001110"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 3713 => y_in <= "10001110"; x_in <= "00000001"; z_correct<="1111111110001110";
        when 3714 => y_in <= "10001110"; x_in <= "00000010"; z_correct<="1111111100011100";
        when 3715 => y_in <= "10001110"; x_in <= "00000011"; z_correct<="1111111010101010";
        when 3716 => y_in <= "10001110"; x_in <= "00000100"; z_correct<="1111111000111000";
        when 3717 => y_in <= "10001110"; x_in <= "00000101"; z_correct<="1111110111000110";
        when 3718 => y_in <= "10001110"; x_in <= "00000110"; z_correct<="1111110101010100";
        when 3719 => y_in <= "10001110"; x_in <= "00000111"; z_correct<="1111110011100010";
        when 3720 => y_in <= "10001110"; x_in <= "00001000"; z_correct<="1111110001110000";
        when 3721 => y_in <= "10001110"; x_in <= "00001001"; z_correct<="1111101111111110";
        when 3722 => y_in <= "10001110"; x_in <= "00001010"; z_correct<="1111101110001100";
        when 3723 => y_in <= "10001110"; x_in <= "00001011"; z_correct<="1111101100011010";
        when 3724 => y_in <= "10001110"; x_in <= "00001100"; z_correct<="1111101010101000";
        when 3725 => y_in <= "10001110"; x_in <= "00001101"; z_correct<="1111101000110110";
        when 3726 => y_in <= "10001110"; x_in <= "00001110"; z_correct<="1111100111000100";
        when 3727 => y_in <= "10001110"; x_in <= "00001111"; z_correct<="1111100101010010";
        when 3728 => y_in <= "10001110"; x_in <= "00010000"; z_correct<="1111100011100000";
        when 3729 => y_in <= "10001110"; x_in <= "00010001"; z_correct<="1111100001101110";
        when 3730 => y_in <= "10001110"; x_in <= "00010010"; z_correct<="1111011111111100";
        when 3731 => y_in <= "10001110"; x_in <= "00010011"; z_correct<="1111011110001010";
        when 3732 => y_in <= "10001110"; x_in <= "00010100"; z_correct<="1111011100011000";
        when 3733 => y_in <= "10001110"; x_in <= "00010101"; z_correct<="1111011010100110";
        when 3734 => y_in <= "10001110"; x_in <= "00010110"; z_correct<="1111011000110100";
        when 3735 => y_in <= "10001110"; x_in <= "00010111"; z_correct<="1111010111000010";
        when 3736 => y_in <= "10001110"; x_in <= "00011000"; z_correct<="1111010101010000";
        when 3737 => y_in <= "10001110"; x_in <= "00011001"; z_correct<="1111010011011110";
        when 3738 => y_in <= "10001110"; x_in <= "00011010"; z_correct<="1111010001101100";
        when 3739 => y_in <= "10001110"; x_in <= "00011011"; z_correct<="1111001111111010";
        when 3740 => y_in <= "10001110"; x_in <= "00011100"; z_correct<="1111001110001000";
        when 3741 => y_in <= "10001110"; x_in <= "00011101"; z_correct<="1111001100010110";
        when 3742 => y_in <= "10001110"; x_in <= "00011110"; z_correct<="1111001010100100";
        when 3743 => y_in <= "10001110"; x_in <= "00011111"; z_correct<="1111001000110010";
        when 3744 => y_in <= "10001110"; x_in <= "00100000"; z_correct<="1111000111000000";
        when 3745 => y_in <= "10001110"; x_in <= "00100001"; z_correct<="1111000101001110";
        when 3746 => y_in <= "10001110"; x_in <= "00100010"; z_correct<="1111000011011100";
        when 3747 => y_in <= "10001110"; x_in <= "00100011"; z_correct<="1111000001101010";
        when 3748 => y_in <= "10001110"; x_in <= "00100100"; z_correct<="1110111111111000";
        when 3749 => y_in <= "10001110"; x_in <= "00100101"; z_correct<="1110111110000110";
        when 3750 => y_in <= "10001110"; x_in <= "00100110"; z_correct<="1110111100010100";
        when 3751 => y_in <= "10001110"; x_in <= "00100111"; z_correct<="1110111010100010";
        when 3752 => y_in <= "10001110"; x_in <= "00101000"; z_correct<="1110111000110000";
        when 3753 => y_in <= "10001110"; x_in <= "00101001"; z_correct<="1110110110111110";
        when 3754 => y_in <= "10001110"; x_in <= "00101010"; z_correct<="1110110101001100";
        when 3755 => y_in <= "10001110"; x_in <= "00101011"; z_correct<="1110110011011010";
        when 3756 => y_in <= "10001110"; x_in <= "00101100"; z_correct<="1110110001101000";
        when 3757 => y_in <= "10001110"; x_in <= "00101101"; z_correct<="1110101111110110";
        when 3758 => y_in <= "10001110"; x_in <= "00101110"; z_correct<="1110101110000100";
        when 3759 => y_in <= "10001110"; x_in <= "00101111"; z_correct<="1110101100010010";
        when 3760 => y_in <= "10001110"; x_in <= "00110000"; z_correct<="1110101010100000";
        when 3761 => y_in <= "10001110"; x_in <= "00110001"; z_correct<="1110101000101110";
        when 3762 => y_in <= "10001110"; x_in <= "00110010"; z_correct<="1110100110111100";
        when 3763 => y_in <= "10001110"; x_in <= "00110011"; z_correct<="1110100101001010";
        when 3764 => y_in <= "10001110"; x_in <= "00110100"; z_correct<="1110100011011000";
        when 3765 => y_in <= "10001110"; x_in <= "00110101"; z_correct<="1110100001100110";
        when 3766 => y_in <= "10001110"; x_in <= "00110110"; z_correct<="1110011111110100";
        when 3767 => y_in <= "10001110"; x_in <= "00110111"; z_correct<="1110011110000010";
        when 3768 => y_in <= "10001110"; x_in <= "00111000"; z_correct<="1110011100010000";
        when 3769 => y_in <= "10001110"; x_in <= "00111001"; z_correct<="1110011010011110";
        when 3770 => y_in <= "10001110"; x_in <= "00111010"; z_correct<="1110011000101100";
        when 3771 => y_in <= "10001110"; x_in <= "00111011"; z_correct<="1110010110111010";
        when 3772 => y_in <= "10001110"; x_in <= "00111100"; z_correct<="1110010101001000";
        when 3773 => y_in <= "10001110"; x_in <= "00111101"; z_correct<="1110010011010110";
        when 3774 => y_in <= "10001110"; x_in <= "00111110"; z_correct<="1110010001100100";
        when 3775 => y_in <= "10001110"; x_in <= "00111111"; z_correct<="1110001111110010";
        when 3776 => y_in <= "10001110"; x_in <= "01000000"; z_correct<="1110001110000000";
        when 3777 => y_in <= "10001110"; x_in <= "01000001"; z_correct<="1110001100001110";
        when 3778 => y_in <= "10001110"; x_in <= "01000010"; z_correct<="1110001010011100";
        when 3779 => y_in <= "10001110"; x_in <= "01000011"; z_correct<="1110001000101010";
        when 3780 => y_in <= "10001110"; x_in <= "01000100"; z_correct<="1110000110111000";
        when 3781 => y_in <= "10001110"; x_in <= "01000101"; z_correct<="1110000101000110";
        when 3782 => y_in <= "10001110"; x_in <= "01000110"; z_correct<="1110000011010100";
        when 3783 => y_in <= "10001110"; x_in <= "01000111"; z_correct<="1110000001100010";
        when 3784 => y_in <= "10001110"; x_in <= "01001000"; z_correct<="1101111111110000";
        when 3785 => y_in <= "10001110"; x_in <= "01001001"; z_correct<="1101111101111110";
        when 3786 => y_in <= "10001110"; x_in <= "01001010"; z_correct<="1101111100001100";
        when 3787 => y_in <= "10001110"; x_in <= "01001011"; z_correct<="1101111010011010";
        when 3788 => y_in <= "10001110"; x_in <= "01001100"; z_correct<="1101111000101000";
        when 3789 => y_in <= "10001110"; x_in <= "01001101"; z_correct<="1101110110110110";
        when 3790 => y_in <= "10001110"; x_in <= "01001110"; z_correct<="1101110101000100";
        when 3791 => y_in <= "10001110"; x_in <= "01001111"; z_correct<="1101110011010010";
        when 3792 => y_in <= "10001110"; x_in <= "01010000"; z_correct<="1101110001100000";
        when 3793 => y_in <= "10001110"; x_in <= "01010001"; z_correct<="1101101111101110";
        when 3794 => y_in <= "10001110"; x_in <= "01010010"; z_correct<="1101101101111100";
        when 3795 => y_in <= "10001110"; x_in <= "01010011"; z_correct<="1101101100001010";
        when 3796 => y_in <= "10001110"; x_in <= "01010100"; z_correct<="1101101010011000";
        when 3797 => y_in <= "10001110"; x_in <= "01010101"; z_correct<="1101101000100110";
        when 3798 => y_in <= "10001110"; x_in <= "01010110"; z_correct<="1101100110110100";
        when 3799 => y_in <= "10001110"; x_in <= "01010111"; z_correct<="1101100101000010";
        when 3800 => y_in <= "10001110"; x_in <= "01011000"; z_correct<="1101100011010000";
        when 3801 => y_in <= "10001110"; x_in <= "01011001"; z_correct<="1101100001011110";
        when 3802 => y_in <= "10001110"; x_in <= "01011010"; z_correct<="1101011111101100";
        when 3803 => y_in <= "10001110"; x_in <= "01011011"; z_correct<="1101011101111010";
        when 3804 => y_in <= "10001110"; x_in <= "01011100"; z_correct<="1101011100001000";
        when 3805 => y_in <= "10001110"; x_in <= "01011101"; z_correct<="1101011010010110";
        when 3806 => y_in <= "10001110"; x_in <= "01011110"; z_correct<="1101011000100100";
        when 3807 => y_in <= "10001110"; x_in <= "01011111"; z_correct<="1101010110110010";
        when 3808 => y_in <= "10001110"; x_in <= "01100000"; z_correct<="1101010101000000";
        when 3809 => y_in <= "10001110"; x_in <= "01100001"; z_correct<="1101010011001110";
        when 3810 => y_in <= "10001110"; x_in <= "01100010"; z_correct<="1101010001011100";
        when 3811 => y_in <= "10001110"; x_in <= "01100011"; z_correct<="1101001111101010";
        when 3812 => y_in <= "10001110"; x_in <= "01100100"; z_correct<="1101001101111000";
        when 3813 => y_in <= "10001110"; x_in <= "01100101"; z_correct<="1101001100000110";
        when 3814 => y_in <= "10001110"; x_in <= "01100110"; z_correct<="1101001010010100";
        when 3815 => y_in <= "10001110"; x_in <= "01100111"; z_correct<="1101001000100010";
        when 3816 => y_in <= "10001110"; x_in <= "01101000"; z_correct<="1101000110110000";
        when 3817 => y_in <= "10001110"; x_in <= "01101001"; z_correct<="1101000100111110";
        when 3818 => y_in <= "10001110"; x_in <= "01101010"; z_correct<="1101000011001100";
        when 3819 => y_in <= "10001110"; x_in <= "01101011"; z_correct<="1101000001011010";
        when 3820 => y_in <= "10001110"; x_in <= "01101100"; z_correct<="1100111111101000";
        when 3821 => y_in <= "10001110"; x_in <= "01101101"; z_correct<="1100111101110110";
        when 3822 => y_in <= "10001110"; x_in <= "01101110"; z_correct<="1100111100000100";
        when 3823 => y_in <= "10001110"; x_in <= "01101111"; z_correct<="1100111010010010";
        when 3824 => y_in <= "10001110"; x_in <= "01110000"; z_correct<="1100111000100000";
        when 3825 => y_in <= "10001110"; x_in <= "01110001"; z_correct<="1100110110101110";
        when 3826 => y_in <= "10001110"; x_in <= "01110010"; z_correct<="1100110100111100";
        when 3827 => y_in <= "10001110"; x_in <= "01110011"; z_correct<="1100110011001010";
        when 3828 => y_in <= "10001110"; x_in <= "01110100"; z_correct<="1100110001011000";
        when 3829 => y_in <= "10001110"; x_in <= "01110101"; z_correct<="1100101111100110";
        when 3830 => y_in <= "10001110"; x_in <= "01110110"; z_correct<="1100101101110100";
        when 3831 => y_in <= "10001110"; x_in <= "01110111"; z_correct<="1100101100000010";
        when 3832 => y_in <= "10001110"; x_in <= "01111000"; z_correct<="1100101010010000";
        when 3833 => y_in <= "10001110"; x_in <= "01111001"; z_correct<="1100101000011110";
        when 3834 => y_in <= "10001110"; x_in <= "01111010"; z_correct<="1100100110101100";
        when 3835 => y_in <= "10001110"; x_in <= "01111011"; z_correct<="1100100100111010";
        when 3836 => y_in <= "10001110"; x_in <= "01111100"; z_correct<="1100100011001000";
        when 3837 => y_in <= "10001110"; x_in <= "01111101"; z_correct<="1100100001010110";
        when 3838 => y_in <= "10001110"; x_in <= "01111110"; z_correct<="1100011111100100";
        when 3839 => y_in <= "10001110"; x_in <= "01111111"; z_correct<="1100011101110010";
        when 3840 => y_in <= "10001111"; x_in <= "10000000"; z_correct<="0011100010000000";
        when 3841 => y_in <= "10001111"; x_in <= "10000001"; z_correct<="0011100000001111";
        when 3842 => y_in <= "10001111"; x_in <= "10000010"; z_correct<="0011011110011110";
        when 3843 => y_in <= "10001111"; x_in <= "10000011"; z_correct<="0011011100101101";
        when 3844 => y_in <= "10001111"; x_in <= "10000100"; z_correct<="0011011010111100";
        when 3845 => y_in <= "10001111"; x_in <= "10000101"; z_correct<="0011011001001011";
        when 3846 => y_in <= "10001111"; x_in <= "10000110"; z_correct<="0011010111011010";
        when 3847 => y_in <= "10001111"; x_in <= "10000111"; z_correct<="0011010101101001";
        when 3848 => y_in <= "10001111"; x_in <= "10001000"; z_correct<="0011010011111000";
        when 3849 => y_in <= "10001111"; x_in <= "10001001"; z_correct<="0011010010000111";
        when 3850 => y_in <= "10001111"; x_in <= "10001010"; z_correct<="0011010000010110";
        when 3851 => y_in <= "10001111"; x_in <= "10001011"; z_correct<="0011001110100101";
        when 3852 => y_in <= "10001111"; x_in <= "10001100"; z_correct<="0011001100110100";
        when 3853 => y_in <= "10001111"; x_in <= "10001101"; z_correct<="0011001011000011";
        when 3854 => y_in <= "10001111"; x_in <= "10001110"; z_correct<="0011001001010010";
        when 3855 => y_in <= "10001111"; x_in <= "10001111"; z_correct<="0011000111100001";
        when 3856 => y_in <= "10001111"; x_in <= "10010000"; z_correct<="0011000101110000";
        when 3857 => y_in <= "10001111"; x_in <= "10010001"; z_correct<="0011000011111111";
        when 3858 => y_in <= "10001111"; x_in <= "10010010"; z_correct<="0011000010001110";
        when 3859 => y_in <= "10001111"; x_in <= "10010011"; z_correct<="0011000000011101";
        when 3860 => y_in <= "10001111"; x_in <= "10010100"; z_correct<="0010111110101100";
        when 3861 => y_in <= "10001111"; x_in <= "10010101"; z_correct<="0010111100111011";
        when 3862 => y_in <= "10001111"; x_in <= "10010110"; z_correct<="0010111011001010";
        when 3863 => y_in <= "10001111"; x_in <= "10010111"; z_correct<="0010111001011001";
        when 3864 => y_in <= "10001111"; x_in <= "10011000"; z_correct<="0010110111101000";
        when 3865 => y_in <= "10001111"; x_in <= "10011001"; z_correct<="0010110101110111";
        when 3866 => y_in <= "10001111"; x_in <= "10011010"; z_correct<="0010110100000110";
        when 3867 => y_in <= "10001111"; x_in <= "10011011"; z_correct<="0010110010010101";
        when 3868 => y_in <= "10001111"; x_in <= "10011100"; z_correct<="0010110000100100";
        when 3869 => y_in <= "10001111"; x_in <= "10011101"; z_correct<="0010101110110011";
        when 3870 => y_in <= "10001111"; x_in <= "10011110"; z_correct<="0010101101000010";
        when 3871 => y_in <= "10001111"; x_in <= "10011111"; z_correct<="0010101011010001";
        when 3872 => y_in <= "10001111"; x_in <= "10100000"; z_correct<="0010101001100000";
        when 3873 => y_in <= "10001111"; x_in <= "10100001"; z_correct<="0010100111101111";
        when 3874 => y_in <= "10001111"; x_in <= "10100010"; z_correct<="0010100101111110";
        when 3875 => y_in <= "10001111"; x_in <= "10100011"; z_correct<="0010100100001101";
        when 3876 => y_in <= "10001111"; x_in <= "10100100"; z_correct<="0010100010011100";
        when 3877 => y_in <= "10001111"; x_in <= "10100101"; z_correct<="0010100000101011";
        when 3878 => y_in <= "10001111"; x_in <= "10100110"; z_correct<="0010011110111010";
        when 3879 => y_in <= "10001111"; x_in <= "10100111"; z_correct<="0010011101001001";
        when 3880 => y_in <= "10001111"; x_in <= "10101000"; z_correct<="0010011011011000";
        when 3881 => y_in <= "10001111"; x_in <= "10101001"; z_correct<="0010011001100111";
        when 3882 => y_in <= "10001111"; x_in <= "10101010"; z_correct<="0010010111110110";
        when 3883 => y_in <= "10001111"; x_in <= "10101011"; z_correct<="0010010110000101";
        when 3884 => y_in <= "10001111"; x_in <= "10101100"; z_correct<="0010010100010100";
        when 3885 => y_in <= "10001111"; x_in <= "10101101"; z_correct<="0010010010100011";
        when 3886 => y_in <= "10001111"; x_in <= "10101110"; z_correct<="0010010000110010";
        when 3887 => y_in <= "10001111"; x_in <= "10101111"; z_correct<="0010001111000001";
        when 3888 => y_in <= "10001111"; x_in <= "10110000"; z_correct<="0010001101010000";
        when 3889 => y_in <= "10001111"; x_in <= "10110001"; z_correct<="0010001011011111";
        when 3890 => y_in <= "10001111"; x_in <= "10110010"; z_correct<="0010001001101110";
        when 3891 => y_in <= "10001111"; x_in <= "10110011"; z_correct<="0010000111111101";
        when 3892 => y_in <= "10001111"; x_in <= "10110100"; z_correct<="0010000110001100";
        when 3893 => y_in <= "10001111"; x_in <= "10110101"; z_correct<="0010000100011011";
        when 3894 => y_in <= "10001111"; x_in <= "10110110"; z_correct<="0010000010101010";
        when 3895 => y_in <= "10001111"; x_in <= "10110111"; z_correct<="0010000000111001";
        when 3896 => y_in <= "10001111"; x_in <= "10111000"; z_correct<="0001111111001000";
        when 3897 => y_in <= "10001111"; x_in <= "10111001"; z_correct<="0001111101010111";
        when 3898 => y_in <= "10001111"; x_in <= "10111010"; z_correct<="0001111011100110";
        when 3899 => y_in <= "10001111"; x_in <= "10111011"; z_correct<="0001111001110101";
        when 3900 => y_in <= "10001111"; x_in <= "10111100"; z_correct<="0001111000000100";
        when 3901 => y_in <= "10001111"; x_in <= "10111101"; z_correct<="0001110110010011";
        when 3902 => y_in <= "10001111"; x_in <= "10111110"; z_correct<="0001110100100010";
        when 3903 => y_in <= "10001111"; x_in <= "10111111"; z_correct<="0001110010110001";
        when 3904 => y_in <= "10001111"; x_in <= "11000000"; z_correct<="0001110001000000";
        when 3905 => y_in <= "10001111"; x_in <= "11000001"; z_correct<="0001101111001111";
        when 3906 => y_in <= "10001111"; x_in <= "11000010"; z_correct<="0001101101011110";
        when 3907 => y_in <= "10001111"; x_in <= "11000011"; z_correct<="0001101011101101";
        when 3908 => y_in <= "10001111"; x_in <= "11000100"; z_correct<="0001101001111100";
        when 3909 => y_in <= "10001111"; x_in <= "11000101"; z_correct<="0001101000001011";
        when 3910 => y_in <= "10001111"; x_in <= "11000110"; z_correct<="0001100110011010";
        when 3911 => y_in <= "10001111"; x_in <= "11000111"; z_correct<="0001100100101001";
        when 3912 => y_in <= "10001111"; x_in <= "11001000"; z_correct<="0001100010111000";
        when 3913 => y_in <= "10001111"; x_in <= "11001001"; z_correct<="0001100001000111";
        when 3914 => y_in <= "10001111"; x_in <= "11001010"; z_correct<="0001011111010110";
        when 3915 => y_in <= "10001111"; x_in <= "11001011"; z_correct<="0001011101100101";
        when 3916 => y_in <= "10001111"; x_in <= "11001100"; z_correct<="0001011011110100";
        when 3917 => y_in <= "10001111"; x_in <= "11001101"; z_correct<="0001011010000011";
        when 3918 => y_in <= "10001111"; x_in <= "11001110"; z_correct<="0001011000010010";
        when 3919 => y_in <= "10001111"; x_in <= "11001111"; z_correct<="0001010110100001";
        when 3920 => y_in <= "10001111"; x_in <= "11010000"; z_correct<="0001010100110000";
        when 3921 => y_in <= "10001111"; x_in <= "11010001"; z_correct<="0001010010111111";
        when 3922 => y_in <= "10001111"; x_in <= "11010010"; z_correct<="0001010001001110";
        when 3923 => y_in <= "10001111"; x_in <= "11010011"; z_correct<="0001001111011101";
        when 3924 => y_in <= "10001111"; x_in <= "11010100"; z_correct<="0001001101101100";
        when 3925 => y_in <= "10001111"; x_in <= "11010101"; z_correct<="0001001011111011";
        when 3926 => y_in <= "10001111"; x_in <= "11010110"; z_correct<="0001001010001010";
        when 3927 => y_in <= "10001111"; x_in <= "11010111"; z_correct<="0001001000011001";
        when 3928 => y_in <= "10001111"; x_in <= "11011000"; z_correct<="0001000110101000";
        when 3929 => y_in <= "10001111"; x_in <= "11011001"; z_correct<="0001000100110111";
        when 3930 => y_in <= "10001111"; x_in <= "11011010"; z_correct<="0001000011000110";
        when 3931 => y_in <= "10001111"; x_in <= "11011011"; z_correct<="0001000001010101";
        when 3932 => y_in <= "10001111"; x_in <= "11011100"; z_correct<="0000111111100100";
        when 3933 => y_in <= "10001111"; x_in <= "11011101"; z_correct<="0000111101110011";
        when 3934 => y_in <= "10001111"; x_in <= "11011110"; z_correct<="0000111100000010";
        when 3935 => y_in <= "10001111"; x_in <= "11011111"; z_correct<="0000111010010001";
        when 3936 => y_in <= "10001111"; x_in <= "11100000"; z_correct<="0000111000100000";
        when 3937 => y_in <= "10001111"; x_in <= "11100001"; z_correct<="0000110110101111";
        when 3938 => y_in <= "10001111"; x_in <= "11100010"; z_correct<="0000110100111110";
        when 3939 => y_in <= "10001111"; x_in <= "11100011"; z_correct<="0000110011001101";
        when 3940 => y_in <= "10001111"; x_in <= "11100100"; z_correct<="0000110001011100";
        when 3941 => y_in <= "10001111"; x_in <= "11100101"; z_correct<="0000101111101011";
        when 3942 => y_in <= "10001111"; x_in <= "11100110"; z_correct<="0000101101111010";
        when 3943 => y_in <= "10001111"; x_in <= "11100111"; z_correct<="0000101100001001";
        when 3944 => y_in <= "10001111"; x_in <= "11101000"; z_correct<="0000101010011000";
        when 3945 => y_in <= "10001111"; x_in <= "11101001"; z_correct<="0000101000100111";
        when 3946 => y_in <= "10001111"; x_in <= "11101010"; z_correct<="0000100110110110";
        when 3947 => y_in <= "10001111"; x_in <= "11101011"; z_correct<="0000100101000101";
        when 3948 => y_in <= "10001111"; x_in <= "11101100"; z_correct<="0000100011010100";
        when 3949 => y_in <= "10001111"; x_in <= "11101101"; z_correct<="0000100001100011";
        when 3950 => y_in <= "10001111"; x_in <= "11101110"; z_correct<="0000011111110010";
        when 3951 => y_in <= "10001111"; x_in <= "11101111"; z_correct<="0000011110000001";
        when 3952 => y_in <= "10001111"; x_in <= "11110000"; z_correct<="0000011100010000";
        when 3953 => y_in <= "10001111"; x_in <= "11110001"; z_correct<="0000011010011111";
        when 3954 => y_in <= "10001111"; x_in <= "11110010"; z_correct<="0000011000101110";
        when 3955 => y_in <= "10001111"; x_in <= "11110011"; z_correct<="0000010110111101";
        when 3956 => y_in <= "10001111"; x_in <= "11110100"; z_correct<="0000010101001100";
        when 3957 => y_in <= "10001111"; x_in <= "11110101"; z_correct<="0000010011011011";
        when 3958 => y_in <= "10001111"; x_in <= "11110110"; z_correct<="0000010001101010";
        when 3959 => y_in <= "10001111"; x_in <= "11110111"; z_correct<="0000001111111001";
        when 3960 => y_in <= "10001111"; x_in <= "11111000"; z_correct<="0000001110001000";
        when 3961 => y_in <= "10001111"; x_in <= "11111001"; z_correct<="0000001100010111";
        when 3962 => y_in <= "10001111"; x_in <= "11111010"; z_correct<="0000001010100110";
        when 3963 => y_in <= "10001111"; x_in <= "11111011"; z_correct<="0000001000110101";
        when 3964 => y_in <= "10001111"; x_in <= "11111100"; z_correct<="0000000111000100";
        when 3965 => y_in <= "10001111"; x_in <= "11111101"; z_correct<="0000000101010011";
        when 3966 => y_in <= "10001111"; x_in <= "11111110"; z_correct<="0000000011100010";
        when 3967 => y_in <= "10001111"; x_in <= "11111111"; z_correct<="0000000001110001";
        when 3968 => y_in <= "10001111"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 3969 => y_in <= "10001111"; x_in <= "00000001"; z_correct<="1111111110001111";
        when 3970 => y_in <= "10001111"; x_in <= "00000010"; z_correct<="1111111100011110";
        when 3971 => y_in <= "10001111"; x_in <= "00000011"; z_correct<="1111111010101101";
        when 3972 => y_in <= "10001111"; x_in <= "00000100"; z_correct<="1111111000111100";
        when 3973 => y_in <= "10001111"; x_in <= "00000101"; z_correct<="1111110111001011";
        when 3974 => y_in <= "10001111"; x_in <= "00000110"; z_correct<="1111110101011010";
        when 3975 => y_in <= "10001111"; x_in <= "00000111"; z_correct<="1111110011101001";
        when 3976 => y_in <= "10001111"; x_in <= "00001000"; z_correct<="1111110001111000";
        when 3977 => y_in <= "10001111"; x_in <= "00001001"; z_correct<="1111110000000111";
        when 3978 => y_in <= "10001111"; x_in <= "00001010"; z_correct<="1111101110010110";
        when 3979 => y_in <= "10001111"; x_in <= "00001011"; z_correct<="1111101100100101";
        when 3980 => y_in <= "10001111"; x_in <= "00001100"; z_correct<="1111101010110100";
        when 3981 => y_in <= "10001111"; x_in <= "00001101"; z_correct<="1111101001000011";
        when 3982 => y_in <= "10001111"; x_in <= "00001110"; z_correct<="1111100111010010";
        when 3983 => y_in <= "10001111"; x_in <= "00001111"; z_correct<="1111100101100001";
        when 3984 => y_in <= "10001111"; x_in <= "00010000"; z_correct<="1111100011110000";
        when 3985 => y_in <= "10001111"; x_in <= "00010001"; z_correct<="1111100001111111";
        when 3986 => y_in <= "10001111"; x_in <= "00010010"; z_correct<="1111100000001110";
        when 3987 => y_in <= "10001111"; x_in <= "00010011"; z_correct<="1111011110011101";
        when 3988 => y_in <= "10001111"; x_in <= "00010100"; z_correct<="1111011100101100";
        when 3989 => y_in <= "10001111"; x_in <= "00010101"; z_correct<="1111011010111011";
        when 3990 => y_in <= "10001111"; x_in <= "00010110"; z_correct<="1111011001001010";
        when 3991 => y_in <= "10001111"; x_in <= "00010111"; z_correct<="1111010111011001";
        when 3992 => y_in <= "10001111"; x_in <= "00011000"; z_correct<="1111010101101000";
        when 3993 => y_in <= "10001111"; x_in <= "00011001"; z_correct<="1111010011110111";
        when 3994 => y_in <= "10001111"; x_in <= "00011010"; z_correct<="1111010010000110";
        when 3995 => y_in <= "10001111"; x_in <= "00011011"; z_correct<="1111010000010101";
        when 3996 => y_in <= "10001111"; x_in <= "00011100"; z_correct<="1111001110100100";
        when 3997 => y_in <= "10001111"; x_in <= "00011101"; z_correct<="1111001100110011";
        when 3998 => y_in <= "10001111"; x_in <= "00011110"; z_correct<="1111001011000010";
        when 3999 => y_in <= "10001111"; x_in <= "00011111"; z_correct<="1111001001010001";
        when 4000 => y_in <= "10001111"; x_in <= "00100000"; z_correct<="1111000111100000";
        when 4001 => y_in <= "10001111"; x_in <= "00100001"; z_correct<="1111000101101111";
        when 4002 => y_in <= "10001111"; x_in <= "00100010"; z_correct<="1111000011111110";
        when 4003 => y_in <= "10001111"; x_in <= "00100011"; z_correct<="1111000010001101";
        when 4004 => y_in <= "10001111"; x_in <= "00100100"; z_correct<="1111000000011100";
        when 4005 => y_in <= "10001111"; x_in <= "00100101"; z_correct<="1110111110101011";
        when 4006 => y_in <= "10001111"; x_in <= "00100110"; z_correct<="1110111100111010";
        when 4007 => y_in <= "10001111"; x_in <= "00100111"; z_correct<="1110111011001001";
        when 4008 => y_in <= "10001111"; x_in <= "00101000"; z_correct<="1110111001011000";
        when 4009 => y_in <= "10001111"; x_in <= "00101001"; z_correct<="1110110111100111";
        when 4010 => y_in <= "10001111"; x_in <= "00101010"; z_correct<="1110110101110110";
        when 4011 => y_in <= "10001111"; x_in <= "00101011"; z_correct<="1110110100000101";
        when 4012 => y_in <= "10001111"; x_in <= "00101100"; z_correct<="1110110010010100";
        when 4013 => y_in <= "10001111"; x_in <= "00101101"; z_correct<="1110110000100011";
        when 4014 => y_in <= "10001111"; x_in <= "00101110"; z_correct<="1110101110110010";
        when 4015 => y_in <= "10001111"; x_in <= "00101111"; z_correct<="1110101101000001";
        when 4016 => y_in <= "10001111"; x_in <= "00110000"; z_correct<="1110101011010000";
        when 4017 => y_in <= "10001111"; x_in <= "00110001"; z_correct<="1110101001011111";
        when 4018 => y_in <= "10001111"; x_in <= "00110010"; z_correct<="1110100111101110";
        when 4019 => y_in <= "10001111"; x_in <= "00110011"; z_correct<="1110100101111101";
        when 4020 => y_in <= "10001111"; x_in <= "00110100"; z_correct<="1110100100001100";
        when 4021 => y_in <= "10001111"; x_in <= "00110101"; z_correct<="1110100010011011";
        when 4022 => y_in <= "10001111"; x_in <= "00110110"; z_correct<="1110100000101010";
        when 4023 => y_in <= "10001111"; x_in <= "00110111"; z_correct<="1110011110111001";
        when 4024 => y_in <= "10001111"; x_in <= "00111000"; z_correct<="1110011101001000";
        when 4025 => y_in <= "10001111"; x_in <= "00111001"; z_correct<="1110011011010111";
        when 4026 => y_in <= "10001111"; x_in <= "00111010"; z_correct<="1110011001100110";
        when 4027 => y_in <= "10001111"; x_in <= "00111011"; z_correct<="1110010111110101";
        when 4028 => y_in <= "10001111"; x_in <= "00111100"; z_correct<="1110010110000100";
        when 4029 => y_in <= "10001111"; x_in <= "00111101"; z_correct<="1110010100010011";
        when 4030 => y_in <= "10001111"; x_in <= "00111110"; z_correct<="1110010010100010";
        when 4031 => y_in <= "10001111"; x_in <= "00111111"; z_correct<="1110010000110001";
        when 4032 => y_in <= "10001111"; x_in <= "01000000"; z_correct<="1110001111000000";
        when 4033 => y_in <= "10001111"; x_in <= "01000001"; z_correct<="1110001101001111";
        when 4034 => y_in <= "10001111"; x_in <= "01000010"; z_correct<="1110001011011110";
        when 4035 => y_in <= "10001111"; x_in <= "01000011"; z_correct<="1110001001101101";
        when 4036 => y_in <= "10001111"; x_in <= "01000100"; z_correct<="1110000111111100";
        when 4037 => y_in <= "10001111"; x_in <= "01000101"; z_correct<="1110000110001011";
        when 4038 => y_in <= "10001111"; x_in <= "01000110"; z_correct<="1110000100011010";
        when 4039 => y_in <= "10001111"; x_in <= "01000111"; z_correct<="1110000010101001";
        when 4040 => y_in <= "10001111"; x_in <= "01001000"; z_correct<="1110000000111000";
        when 4041 => y_in <= "10001111"; x_in <= "01001001"; z_correct<="1101111111000111";
        when 4042 => y_in <= "10001111"; x_in <= "01001010"; z_correct<="1101111101010110";
        when 4043 => y_in <= "10001111"; x_in <= "01001011"; z_correct<="1101111011100101";
        when 4044 => y_in <= "10001111"; x_in <= "01001100"; z_correct<="1101111001110100";
        when 4045 => y_in <= "10001111"; x_in <= "01001101"; z_correct<="1101111000000011";
        when 4046 => y_in <= "10001111"; x_in <= "01001110"; z_correct<="1101110110010010";
        when 4047 => y_in <= "10001111"; x_in <= "01001111"; z_correct<="1101110100100001";
        when 4048 => y_in <= "10001111"; x_in <= "01010000"; z_correct<="1101110010110000";
        when 4049 => y_in <= "10001111"; x_in <= "01010001"; z_correct<="1101110000111111";
        when 4050 => y_in <= "10001111"; x_in <= "01010010"; z_correct<="1101101111001110";
        when 4051 => y_in <= "10001111"; x_in <= "01010011"; z_correct<="1101101101011101";
        when 4052 => y_in <= "10001111"; x_in <= "01010100"; z_correct<="1101101011101100";
        when 4053 => y_in <= "10001111"; x_in <= "01010101"; z_correct<="1101101001111011";
        when 4054 => y_in <= "10001111"; x_in <= "01010110"; z_correct<="1101101000001010";
        when 4055 => y_in <= "10001111"; x_in <= "01010111"; z_correct<="1101100110011001";
        when 4056 => y_in <= "10001111"; x_in <= "01011000"; z_correct<="1101100100101000";
        when 4057 => y_in <= "10001111"; x_in <= "01011001"; z_correct<="1101100010110111";
        when 4058 => y_in <= "10001111"; x_in <= "01011010"; z_correct<="1101100001000110";
        when 4059 => y_in <= "10001111"; x_in <= "01011011"; z_correct<="1101011111010101";
        when 4060 => y_in <= "10001111"; x_in <= "01011100"; z_correct<="1101011101100100";
        when 4061 => y_in <= "10001111"; x_in <= "01011101"; z_correct<="1101011011110011";
        when 4062 => y_in <= "10001111"; x_in <= "01011110"; z_correct<="1101011010000010";
        when 4063 => y_in <= "10001111"; x_in <= "01011111"; z_correct<="1101011000010001";
        when 4064 => y_in <= "10001111"; x_in <= "01100000"; z_correct<="1101010110100000";
        when 4065 => y_in <= "10001111"; x_in <= "01100001"; z_correct<="1101010100101111";
        when 4066 => y_in <= "10001111"; x_in <= "01100010"; z_correct<="1101010010111110";
        when 4067 => y_in <= "10001111"; x_in <= "01100011"; z_correct<="1101010001001101";
        when 4068 => y_in <= "10001111"; x_in <= "01100100"; z_correct<="1101001111011100";
        when 4069 => y_in <= "10001111"; x_in <= "01100101"; z_correct<="1101001101101011";
        when 4070 => y_in <= "10001111"; x_in <= "01100110"; z_correct<="1101001011111010";
        when 4071 => y_in <= "10001111"; x_in <= "01100111"; z_correct<="1101001010001001";
        when 4072 => y_in <= "10001111"; x_in <= "01101000"; z_correct<="1101001000011000";
        when 4073 => y_in <= "10001111"; x_in <= "01101001"; z_correct<="1101000110100111";
        when 4074 => y_in <= "10001111"; x_in <= "01101010"; z_correct<="1101000100110110";
        when 4075 => y_in <= "10001111"; x_in <= "01101011"; z_correct<="1101000011000101";
        when 4076 => y_in <= "10001111"; x_in <= "01101100"; z_correct<="1101000001010100";
        when 4077 => y_in <= "10001111"; x_in <= "01101101"; z_correct<="1100111111100011";
        when 4078 => y_in <= "10001111"; x_in <= "01101110"; z_correct<="1100111101110010";
        when 4079 => y_in <= "10001111"; x_in <= "01101111"; z_correct<="1100111100000001";
        when 4080 => y_in <= "10001111"; x_in <= "01110000"; z_correct<="1100111010010000";
        when 4081 => y_in <= "10001111"; x_in <= "01110001"; z_correct<="1100111000011111";
        when 4082 => y_in <= "10001111"; x_in <= "01110010"; z_correct<="1100110110101110";
        when 4083 => y_in <= "10001111"; x_in <= "01110011"; z_correct<="1100110100111101";
        when 4084 => y_in <= "10001111"; x_in <= "01110100"; z_correct<="1100110011001100";
        when 4085 => y_in <= "10001111"; x_in <= "01110101"; z_correct<="1100110001011011";
        when 4086 => y_in <= "10001111"; x_in <= "01110110"; z_correct<="1100101111101010";
        when 4087 => y_in <= "10001111"; x_in <= "01110111"; z_correct<="1100101101111001";
        when 4088 => y_in <= "10001111"; x_in <= "01111000"; z_correct<="1100101100001000";
        when 4089 => y_in <= "10001111"; x_in <= "01111001"; z_correct<="1100101010010111";
        when 4090 => y_in <= "10001111"; x_in <= "01111010"; z_correct<="1100101000100110";
        when 4091 => y_in <= "10001111"; x_in <= "01111011"; z_correct<="1100100110110101";
        when 4092 => y_in <= "10001111"; x_in <= "01111100"; z_correct<="1100100101000100";
        when 4093 => y_in <= "10001111"; x_in <= "01111101"; z_correct<="1100100011010011";
        when 4094 => y_in <= "10001111"; x_in <= "01111110"; z_correct<="1100100001100010";
        when 4095 => y_in <= "10001111"; x_in <= "01111111"; z_correct<="1100011111110001";
        when 4096 => y_in <= "10010000"; x_in <= "10000000"; z_correct<="0011100000000000";
        when 4097 => y_in <= "10010000"; x_in <= "10000001"; z_correct<="0011011110010000";
        when 4098 => y_in <= "10010000"; x_in <= "10000010"; z_correct<="0011011100100000";
        when 4099 => y_in <= "10010000"; x_in <= "10000011"; z_correct<="0011011010110000";
        when 4100 => y_in <= "10010000"; x_in <= "10000100"; z_correct<="0011011001000000";
        when 4101 => y_in <= "10010000"; x_in <= "10000101"; z_correct<="0011010111010000";
        when 4102 => y_in <= "10010000"; x_in <= "10000110"; z_correct<="0011010101100000";
        when 4103 => y_in <= "10010000"; x_in <= "10000111"; z_correct<="0011010011110000";
        when 4104 => y_in <= "10010000"; x_in <= "10001000"; z_correct<="0011010010000000";
        when 4105 => y_in <= "10010000"; x_in <= "10001001"; z_correct<="0011010000010000";
        when 4106 => y_in <= "10010000"; x_in <= "10001010"; z_correct<="0011001110100000";
        when 4107 => y_in <= "10010000"; x_in <= "10001011"; z_correct<="0011001100110000";
        when 4108 => y_in <= "10010000"; x_in <= "10001100"; z_correct<="0011001011000000";
        when 4109 => y_in <= "10010000"; x_in <= "10001101"; z_correct<="0011001001010000";
        when 4110 => y_in <= "10010000"; x_in <= "10001110"; z_correct<="0011000111100000";
        when 4111 => y_in <= "10010000"; x_in <= "10001111"; z_correct<="0011000101110000";
        when 4112 => y_in <= "10010000"; x_in <= "10010000"; z_correct<="0011000100000000";
        when 4113 => y_in <= "10010000"; x_in <= "10010001"; z_correct<="0011000010010000";
        when 4114 => y_in <= "10010000"; x_in <= "10010010"; z_correct<="0011000000100000";
        when 4115 => y_in <= "10010000"; x_in <= "10010011"; z_correct<="0010111110110000";
        when 4116 => y_in <= "10010000"; x_in <= "10010100"; z_correct<="0010111101000000";
        when 4117 => y_in <= "10010000"; x_in <= "10010101"; z_correct<="0010111011010000";
        when 4118 => y_in <= "10010000"; x_in <= "10010110"; z_correct<="0010111001100000";
        when 4119 => y_in <= "10010000"; x_in <= "10010111"; z_correct<="0010110111110000";
        when 4120 => y_in <= "10010000"; x_in <= "10011000"; z_correct<="0010110110000000";
        when 4121 => y_in <= "10010000"; x_in <= "10011001"; z_correct<="0010110100010000";
        when 4122 => y_in <= "10010000"; x_in <= "10011010"; z_correct<="0010110010100000";
        when 4123 => y_in <= "10010000"; x_in <= "10011011"; z_correct<="0010110000110000";
        when 4124 => y_in <= "10010000"; x_in <= "10011100"; z_correct<="0010101111000000";
        when 4125 => y_in <= "10010000"; x_in <= "10011101"; z_correct<="0010101101010000";
        when 4126 => y_in <= "10010000"; x_in <= "10011110"; z_correct<="0010101011100000";
        when 4127 => y_in <= "10010000"; x_in <= "10011111"; z_correct<="0010101001110000";
        when 4128 => y_in <= "10010000"; x_in <= "10100000"; z_correct<="0010101000000000";
        when 4129 => y_in <= "10010000"; x_in <= "10100001"; z_correct<="0010100110010000";
        when 4130 => y_in <= "10010000"; x_in <= "10100010"; z_correct<="0010100100100000";
        when 4131 => y_in <= "10010000"; x_in <= "10100011"; z_correct<="0010100010110000";
        when 4132 => y_in <= "10010000"; x_in <= "10100100"; z_correct<="0010100001000000";
        when 4133 => y_in <= "10010000"; x_in <= "10100101"; z_correct<="0010011111010000";
        when 4134 => y_in <= "10010000"; x_in <= "10100110"; z_correct<="0010011101100000";
        when 4135 => y_in <= "10010000"; x_in <= "10100111"; z_correct<="0010011011110000";
        when 4136 => y_in <= "10010000"; x_in <= "10101000"; z_correct<="0010011010000000";
        when 4137 => y_in <= "10010000"; x_in <= "10101001"; z_correct<="0010011000010000";
        when 4138 => y_in <= "10010000"; x_in <= "10101010"; z_correct<="0010010110100000";
        when 4139 => y_in <= "10010000"; x_in <= "10101011"; z_correct<="0010010100110000";
        when 4140 => y_in <= "10010000"; x_in <= "10101100"; z_correct<="0010010011000000";
        when 4141 => y_in <= "10010000"; x_in <= "10101101"; z_correct<="0010010001010000";
        when 4142 => y_in <= "10010000"; x_in <= "10101110"; z_correct<="0010001111100000";
        when 4143 => y_in <= "10010000"; x_in <= "10101111"; z_correct<="0010001101110000";
        when 4144 => y_in <= "10010000"; x_in <= "10110000"; z_correct<="0010001100000000";
        when 4145 => y_in <= "10010000"; x_in <= "10110001"; z_correct<="0010001010010000";
        when 4146 => y_in <= "10010000"; x_in <= "10110010"; z_correct<="0010001000100000";
        when 4147 => y_in <= "10010000"; x_in <= "10110011"; z_correct<="0010000110110000";
        when 4148 => y_in <= "10010000"; x_in <= "10110100"; z_correct<="0010000101000000";
        when 4149 => y_in <= "10010000"; x_in <= "10110101"; z_correct<="0010000011010000";
        when 4150 => y_in <= "10010000"; x_in <= "10110110"; z_correct<="0010000001100000";
        when 4151 => y_in <= "10010000"; x_in <= "10110111"; z_correct<="0001111111110000";
        when 4152 => y_in <= "10010000"; x_in <= "10111000"; z_correct<="0001111110000000";
        when 4153 => y_in <= "10010000"; x_in <= "10111001"; z_correct<="0001111100010000";
        when 4154 => y_in <= "10010000"; x_in <= "10111010"; z_correct<="0001111010100000";
        when 4155 => y_in <= "10010000"; x_in <= "10111011"; z_correct<="0001111000110000";
        when 4156 => y_in <= "10010000"; x_in <= "10111100"; z_correct<="0001110111000000";
        when 4157 => y_in <= "10010000"; x_in <= "10111101"; z_correct<="0001110101010000";
        when 4158 => y_in <= "10010000"; x_in <= "10111110"; z_correct<="0001110011100000";
        when 4159 => y_in <= "10010000"; x_in <= "10111111"; z_correct<="0001110001110000";
        when 4160 => y_in <= "10010000"; x_in <= "11000000"; z_correct<="0001110000000000";
        when 4161 => y_in <= "10010000"; x_in <= "11000001"; z_correct<="0001101110010000";
        when 4162 => y_in <= "10010000"; x_in <= "11000010"; z_correct<="0001101100100000";
        when 4163 => y_in <= "10010000"; x_in <= "11000011"; z_correct<="0001101010110000";
        when 4164 => y_in <= "10010000"; x_in <= "11000100"; z_correct<="0001101001000000";
        when 4165 => y_in <= "10010000"; x_in <= "11000101"; z_correct<="0001100111010000";
        when 4166 => y_in <= "10010000"; x_in <= "11000110"; z_correct<="0001100101100000";
        when 4167 => y_in <= "10010000"; x_in <= "11000111"; z_correct<="0001100011110000";
        when 4168 => y_in <= "10010000"; x_in <= "11001000"; z_correct<="0001100010000000";
        when 4169 => y_in <= "10010000"; x_in <= "11001001"; z_correct<="0001100000010000";
        when 4170 => y_in <= "10010000"; x_in <= "11001010"; z_correct<="0001011110100000";
        when 4171 => y_in <= "10010000"; x_in <= "11001011"; z_correct<="0001011100110000";
        when 4172 => y_in <= "10010000"; x_in <= "11001100"; z_correct<="0001011011000000";
        when 4173 => y_in <= "10010000"; x_in <= "11001101"; z_correct<="0001011001010000";
        when 4174 => y_in <= "10010000"; x_in <= "11001110"; z_correct<="0001010111100000";
        when 4175 => y_in <= "10010000"; x_in <= "11001111"; z_correct<="0001010101110000";
        when 4176 => y_in <= "10010000"; x_in <= "11010000"; z_correct<="0001010100000000";
        when 4177 => y_in <= "10010000"; x_in <= "11010001"; z_correct<="0001010010010000";
        when 4178 => y_in <= "10010000"; x_in <= "11010010"; z_correct<="0001010000100000";
        when 4179 => y_in <= "10010000"; x_in <= "11010011"; z_correct<="0001001110110000";
        when 4180 => y_in <= "10010000"; x_in <= "11010100"; z_correct<="0001001101000000";
        when 4181 => y_in <= "10010000"; x_in <= "11010101"; z_correct<="0001001011010000";
        when 4182 => y_in <= "10010000"; x_in <= "11010110"; z_correct<="0001001001100000";
        when 4183 => y_in <= "10010000"; x_in <= "11010111"; z_correct<="0001000111110000";
        when 4184 => y_in <= "10010000"; x_in <= "11011000"; z_correct<="0001000110000000";
        when 4185 => y_in <= "10010000"; x_in <= "11011001"; z_correct<="0001000100010000";
        when 4186 => y_in <= "10010000"; x_in <= "11011010"; z_correct<="0001000010100000";
        when 4187 => y_in <= "10010000"; x_in <= "11011011"; z_correct<="0001000000110000";
        when 4188 => y_in <= "10010000"; x_in <= "11011100"; z_correct<="0000111111000000";
        when 4189 => y_in <= "10010000"; x_in <= "11011101"; z_correct<="0000111101010000";
        when 4190 => y_in <= "10010000"; x_in <= "11011110"; z_correct<="0000111011100000";
        when 4191 => y_in <= "10010000"; x_in <= "11011111"; z_correct<="0000111001110000";
        when 4192 => y_in <= "10010000"; x_in <= "11100000"; z_correct<="0000111000000000";
        when 4193 => y_in <= "10010000"; x_in <= "11100001"; z_correct<="0000110110010000";
        when 4194 => y_in <= "10010000"; x_in <= "11100010"; z_correct<="0000110100100000";
        when 4195 => y_in <= "10010000"; x_in <= "11100011"; z_correct<="0000110010110000";
        when 4196 => y_in <= "10010000"; x_in <= "11100100"; z_correct<="0000110001000000";
        when 4197 => y_in <= "10010000"; x_in <= "11100101"; z_correct<="0000101111010000";
        when 4198 => y_in <= "10010000"; x_in <= "11100110"; z_correct<="0000101101100000";
        when 4199 => y_in <= "10010000"; x_in <= "11100111"; z_correct<="0000101011110000";
        when 4200 => y_in <= "10010000"; x_in <= "11101000"; z_correct<="0000101010000000";
        when 4201 => y_in <= "10010000"; x_in <= "11101001"; z_correct<="0000101000010000";
        when 4202 => y_in <= "10010000"; x_in <= "11101010"; z_correct<="0000100110100000";
        when 4203 => y_in <= "10010000"; x_in <= "11101011"; z_correct<="0000100100110000";
        when 4204 => y_in <= "10010000"; x_in <= "11101100"; z_correct<="0000100011000000";
        when 4205 => y_in <= "10010000"; x_in <= "11101101"; z_correct<="0000100001010000";
        when 4206 => y_in <= "10010000"; x_in <= "11101110"; z_correct<="0000011111100000";
        when 4207 => y_in <= "10010000"; x_in <= "11101111"; z_correct<="0000011101110000";
        when 4208 => y_in <= "10010000"; x_in <= "11110000"; z_correct<="0000011100000000";
        when 4209 => y_in <= "10010000"; x_in <= "11110001"; z_correct<="0000011010010000";
        when 4210 => y_in <= "10010000"; x_in <= "11110010"; z_correct<="0000011000100000";
        when 4211 => y_in <= "10010000"; x_in <= "11110011"; z_correct<="0000010110110000";
        when 4212 => y_in <= "10010000"; x_in <= "11110100"; z_correct<="0000010101000000";
        when 4213 => y_in <= "10010000"; x_in <= "11110101"; z_correct<="0000010011010000";
        when 4214 => y_in <= "10010000"; x_in <= "11110110"; z_correct<="0000010001100000";
        when 4215 => y_in <= "10010000"; x_in <= "11110111"; z_correct<="0000001111110000";
        when 4216 => y_in <= "10010000"; x_in <= "11111000"; z_correct<="0000001110000000";
        when 4217 => y_in <= "10010000"; x_in <= "11111001"; z_correct<="0000001100010000";
        when 4218 => y_in <= "10010000"; x_in <= "11111010"; z_correct<="0000001010100000";
        when 4219 => y_in <= "10010000"; x_in <= "11111011"; z_correct<="0000001000110000";
        when 4220 => y_in <= "10010000"; x_in <= "11111100"; z_correct<="0000000111000000";
        when 4221 => y_in <= "10010000"; x_in <= "11111101"; z_correct<="0000000101010000";
        when 4222 => y_in <= "10010000"; x_in <= "11111110"; z_correct<="0000000011100000";
        when 4223 => y_in <= "10010000"; x_in <= "11111111"; z_correct<="0000000001110000";
        when 4224 => y_in <= "10010000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 4225 => y_in <= "10010000"; x_in <= "00000001"; z_correct<="1111111110010000";
        when 4226 => y_in <= "10010000"; x_in <= "00000010"; z_correct<="1111111100100000";
        when 4227 => y_in <= "10010000"; x_in <= "00000011"; z_correct<="1111111010110000";
        when 4228 => y_in <= "10010000"; x_in <= "00000100"; z_correct<="1111111001000000";
        when 4229 => y_in <= "10010000"; x_in <= "00000101"; z_correct<="1111110111010000";
        when 4230 => y_in <= "10010000"; x_in <= "00000110"; z_correct<="1111110101100000";
        when 4231 => y_in <= "10010000"; x_in <= "00000111"; z_correct<="1111110011110000";
        when 4232 => y_in <= "10010000"; x_in <= "00001000"; z_correct<="1111110010000000";
        when 4233 => y_in <= "10010000"; x_in <= "00001001"; z_correct<="1111110000010000";
        when 4234 => y_in <= "10010000"; x_in <= "00001010"; z_correct<="1111101110100000";
        when 4235 => y_in <= "10010000"; x_in <= "00001011"; z_correct<="1111101100110000";
        when 4236 => y_in <= "10010000"; x_in <= "00001100"; z_correct<="1111101011000000";
        when 4237 => y_in <= "10010000"; x_in <= "00001101"; z_correct<="1111101001010000";
        when 4238 => y_in <= "10010000"; x_in <= "00001110"; z_correct<="1111100111100000";
        when 4239 => y_in <= "10010000"; x_in <= "00001111"; z_correct<="1111100101110000";
        when 4240 => y_in <= "10010000"; x_in <= "00010000"; z_correct<="1111100100000000";
        when 4241 => y_in <= "10010000"; x_in <= "00010001"; z_correct<="1111100010010000";
        when 4242 => y_in <= "10010000"; x_in <= "00010010"; z_correct<="1111100000100000";
        when 4243 => y_in <= "10010000"; x_in <= "00010011"; z_correct<="1111011110110000";
        when 4244 => y_in <= "10010000"; x_in <= "00010100"; z_correct<="1111011101000000";
        when 4245 => y_in <= "10010000"; x_in <= "00010101"; z_correct<="1111011011010000";
        when 4246 => y_in <= "10010000"; x_in <= "00010110"; z_correct<="1111011001100000";
        when 4247 => y_in <= "10010000"; x_in <= "00010111"; z_correct<="1111010111110000";
        when 4248 => y_in <= "10010000"; x_in <= "00011000"; z_correct<="1111010110000000";
        when 4249 => y_in <= "10010000"; x_in <= "00011001"; z_correct<="1111010100010000";
        when 4250 => y_in <= "10010000"; x_in <= "00011010"; z_correct<="1111010010100000";
        when 4251 => y_in <= "10010000"; x_in <= "00011011"; z_correct<="1111010000110000";
        when 4252 => y_in <= "10010000"; x_in <= "00011100"; z_correct<="1111001111000000";
        when 4253 => y_in <= "10010000"; x_in <= "00011101"; z_correct<="1111001101010000";
        when 4254 => y_in <= "10010000"; x_in <= "00011110"; z_correct<="1111001011100000";
        when 4255 => y_in <= "10010000"; x_in <= "00011111"; z_correct<="1111001001110000";
        when 4256 => y_in <= "10010000"; x_in <= "00100000"; z_correct<="1111001000000000";
        when 4257 => y_in <= "10010000"; x_in <= "00100001"; z_correct<="1111000110010000";
        when 4258 => y_in <= "10010000"; x_in <= "00100010"; z_correct<="1111000100100000";
        when 4259 => y_in <= "10010000"; x_in <= "00100011"; z_correct<="1111000010110000";
        when 4260 => y_in <= "10010000"; x_in <= "00100100"; z_correct<="1111000001000000";
        when 4261 => y_in <= "10010000"; x_in <= "00100101"; z_correct<="1110111111010000";
        when 4262 => y_in <= "10010000"; x_in <= "00100110"; z_correct<="1110111101100000";
        when 4263 => y_in <= "10010000"; x_in <= "00100111"; z_correct<="1110111011110000";
        when 4264 => y_in <= "10010000"; x_in <= "00101000"; z_correct<="1110111010000000";
        when 4265 => y_in <= "10010000"; x_in <= "00101001"; z_correct<="1110111000010000";
        when 4266 => y_in <= "10010000"; x_in <= "00101010"; z_correct<="1110110110100000";
        when 4267 => y_in <= "10010000"; x_in <= "00101011"; z_correct<="1110110100110000";
        when 4268 => y_in <= "10010000"; x_in <= "00101100"; z_correct<="1110110011000000";
        when 4269 => y_in <= "10010000"; x_in <= "00101101"; z_correct<="1110110001010000";
        when 4270 => y_in <= "10010000"; x_in <= "00101110"; z_correct<="1110101111100000";
        when 4271 => y_in <= "10010000"; x_in <= "00101111"; z_correct<="1110101101110000";
        when 4272 => y_in <= "10010000"; x_in <= "00110000"; z_correct<="1110101100000000";
        when 4273 => y_in <= "10010000"; x_in <= "00110001"; z_correct<="1110101010010000";
        when 4274 => y_in <= "10010000"; x_in <= "00110010"; z_correct<="1110101000100000";
        when 4275 => y_in <= "10010000"; x_in <= "00110011"; z_correct<="1110100110110000";
        when 4276 => y_in <= "10010000"; x_in <= "00110100"; z_correct<="1110100101000000";
        when 4277 => y_in <= "10010000"; x_in <= "00110101"; z_correct<="1110100011010000";
        when 4278 => y_in <= "10010000"; x_in <= "00110110"; z_correct<="1110100001100000";
        when 4279 => y_in <= "10010000"; x_in <= "00110111"; z_correct<="1110011111110000";
        when 4280 => y_in <= "10010000"; x_in <= "00111000"; z_correct<="1110011110000000";
        when 4281 => y_in <= "10010000"; x_in <= "00111001"; z_correct<="1110011100010000";
        when 4282 => y_in <= "10010000"; x_in <= "00111010"; z_correct<="1110011010100000";
        when 4283 => y_in <= "10010000"; x_in <= "00111011"; z_correct<="1110011000110000";
        when 4284 => y_in <= "10010000"; x_in <= "00111100"; z_correct<="1110010111000000";
        when 4285 => y_in <= "10010000"; x_in <= "00111101"; z_correct<="1110010101010000";
        when 4286 => y_in <= "10010000"; x_in <= "00111110"; z_correct<="1110010011100000";
        when 4287 => y_in <= "10010000"; x_in <= "00111111"; z_correct<="1110010001110000";
        when 4288 => y_in <= "10010000"; x_in <= "01000000"; z_correct<="1110010000000000";
        when 4289 => y_in <= "10010000"; x_in <= "01000001"; z_correct<="1110001110010000";
        when 4290 => y_in <= "10010000"; x_in <= "01000010"; z_correct<="1110001100100000";
        when 4291 => y_in <= "10010000"; x_in <= "01000011"; z_correct<="1110001010110000";
        when 4292 => y_in <= "10010000"; x_in <= "01000100"; z_correct<="1110001001000000";
        when 4293 => y_in <= "10010000"; x_in <= "01000101"; z_correct<="1110000111010000";
        when 4294 => y_in <= "10010000"; x_in <= "01000110"; z_correct<="1110000101100000";
        when 4295 => y_in <= "10010000"; x_in <= "01000111"; z_correct<="1110000011110000";
        when 4296 => y_in <= "10010000"; x_in <= "01001000"; z_correct<="1110000010000000";
        when 4297 => y_in <= "10010000"; x_in <= "01001001"; z_correct<="1110000000010000";
        when 4298 => y_in <= "10010000"; x_in <= "01001010"; z_correct<="1101111110100000";
        when 4299 => y_in <= "10010000"; x_in <= "01001011"; z_correct<="1101111100110000";
        when 4300 => y_in <= "10010000"; x_in <= "01001100"; z_correct<="1101111011000000";
        when 4301 => y_in <= "10010000"; x_in <= "01001101"; z_correct<="1101111001010000";
        when 4302 => y_in <= "10010000"; x_in <= "01001110"; z_correct<="1101110111100000";
        when 4303 => y_in <= "10010000"; x_in <= "01001111"; z_correct<="1101110101110000";
        when 4304 => y_in <= "10010000"; x_in <= "01010000"; z_correct<="1101110100000000";
        when 4305 => y_in <= "10010000"; x_in <= "01010001"; z_correct<="1101110010010000";
        when 4306 => y_in <= "10010000"; x_in <= "01010010"; z_correct<="1101110000100000";
        when 4307 => y_in <= "10010000"; x_in <= "01010011"; z_correct<="1101101110110000";
        when 4308 => y_in <= "10010000"; x_in <= "01010100"; z_correct<="1101101101000000";
        when 4309 => y_in <= "10010000"; x_in <= "01010101"; z_correct<="1101101011010000";
        when 4310 => y_in <= "10010000"; x_in <= "01010110"; z_correct<="1101101001100000";
        when 4311 => y_in <= "10010000"; x_in <= "01010111"; z_correct<="1101100111110000";
        when 4312 => y_in <= "10010000"; x_in <= "01011000"; z_correct<="1101100110000000";
        when 4313 => y_in <= "10010000"; x_in <= "01011001"; z_correct<="1101100100010000";
        when 4314 => y_in <= "10010000"; x_in <= "01011010"; z_correct<="1101100010100000";
        when 4315 => y_in <= "10010000"; x_in <= "01011011"; z_correct<="1101100000110000";
        when 4316 => y_in <= "10010000"; x_in <= "01011100"; z_correct<="1101011111000000";
        when 4317 => y_in <= "10010000"; x_in <= "01011101"; z_correct<="1101011101010000";
        when 4318 => y_in <= "10010000"; x_in <= "01011110"; z_correct<="1101011011100000";
        when 4319 => y_in <= "10010000"; x_in <= "01011111"; z_correct<="1101011001110000";
        when 4320 => y_in <= "10010000"; x_in <= "01100000"; z_correct<="1101011000000000";
        when 4321 => y_in <= "10010000"; x_in <= "01100001"; z_correct<="1101010110010000";
        when 4322 => y_in <= "10010000"; x_in <= "01100010"; z_correct<="1101010100100000";
        when 4323 => y_in <= "10010000"; x_in <= "01100011"; z_correct<="1101010010110000";
        when 4324 => y_in <= "10010000"; x_in <= "01100100"; z_correct<="1101010001000000";
        when 4325 => y_in <= "10010000"; x_in <= "01100101"; z_correct<="1101001111010000";
        when 4326 => y_in <= "10010000"; x_in <= "01100110"; z_correct<="1101001101100000";
        when 4327 => y_in <= "10010000"; x_in <= "01100111"; z_correct<="1101001011110000";
        when 4328 => y_in <= "10010000"; x_in <= "01101000"; z_correct<="1101001010000000";
        when 4329 => y_in <= "10010000"; x_in <= "01101001"; z_correct<="1101001000010000";
        when 4330 => y_in <= "10010000"; x_in <= "01101010"; z_correct<="1101000110100000";
        when 4331 => y_in <= "10010000"; x_in <= "01101011"; z_correct<="1101000100110000";
        when 4332 => y_in <= "10010000"; x_in <= "01101100"; z_correct<="1101000011000000";
        when 4333 => y_in <= "10010000"; x_in <= "01101101"; z_correct<="1101000001010000";
        when 4334 => y_in <= "10010000"; x_in <= "01101110"; z_correct<="1100111111100000";
        when 4335 => y_in <= "10010000"; x_in <= "01101111"; z_correct<="1100111101110000";
        when 4336 => y_in <= "10010000"; x_in <= "01110000"; z_correct<="1100111100000000";
        when 4337 => y_in <= "10010000"; x_in <= "01110001"; z_correct<="1100111010010000";
        when 4338 => y_in <= "10010000"; x_in <= "01110010"; z_correct<="1100111000100000";
        when 4339 => y_in <= "10010000"; x_in <= "01110011"; z_correct<="1100110110110000";
        when 4340 => y_in <= "10010000"; x_in <= "01110100"; z_correct<="1100110101000000";
        when 4341 => y_in <= "10010000"; x_in <= "01110101"; z_correct<="1100110011010000";
        when 4342 => y_in <= "10010000"; x_in <= "01110110"; z_correct<="1100110001100000";
        when 4343 => y_in <= "10010000"; x_in <= "01110111"; z_correct<="1100101111110000";
        when 4344 => y_in <= "10010000"; x_in <= "01111000"; z_correct<="1100101110000000";
        when 4345 => y_in <= "10010000"; x_in <= "01111001"; z_correct<="1100101100010000";
        when 4346 => y_in <= "10010000"; x_in <= "01111010"; z_correct<="1100101010100000";
        when 4347 => y_in <= "10010000"; x_in <= "01111011"; z_correct<="1100101000110000";
        when 4348 => y_in <= "10010000"; x_in <= "01111100"; z_correct<="1100100111000000";
        when 4349 => y_in <= "10010000"; x_in <= "01111101"; z_correct<="1100100101010000";
        when 4350 => y_in <= "10010000"; x_in <= "01111110"; z_correct<="1100100011100000";
        when 4351 => y_in <= "10010000"; x_in <= "01111111"; z_correct<="1100100001110000";
        when 4352 => y_in <= "10010001"; x_in <= "10000000"; z_correct<="0011011110000000";
        when 4353 => y_in <= "10010001"; x_in <= "10000001"; z_correct<="0011011100010001";
        when 4354 => y_in <= "10010001"; x_in <= "10000010"; z_correct<="0011011010100010";
        when 4355 => y_in <= "10010001"; x_in <= "10000011"; z_correct<="0011011000110011";
        when 4356 => y_in <= "10010001"; x_in <= "10000100"; z_correct<="0011010111000100";
        when 4357 => y_in <= "10010001"; x_in <= "10000101"; z_correct<="0011010101010101";
        when 4358 => y_in <= "10010001"; x_in <= "10000110"; z_correct<="0011010011100110";
        when 4359 => y_in <= "10010001"; x_in <= "10000111"; z_correct<="0011010001110111";
        when 4360 => y_in <= "10010001"; x_in <= "10001000"; z_correct<="0011010000001000";
        when 4361 => y_in <= "10010001"; x_in <= "10001001"; z_correct<="0011001110011001";
        when 4362 => y_in <= "10010001"; x_in <= "10001010"; z_correct<="0011001100101010";
        when 4363 => y_in <= "10010001"; x_in <= "10001011"; z_correct<="0011001010111011";
        when 4364 => y_in <= "10010001"; x_in <= "10001100"; z_correct<="0011001001001100";
        when 4365 => y_in <= "10010001"; x_in <= "10001101"; z_correct<="0011000111011101";
        when 4366 => y_in <= "10010001"; x_in <= "10001110"; z_correct<="0011000101101110";
        when 4367 => y_in <= "10010001"; x_in <= "10001111"; z_correct<="0011000011111111";
        when 4368 => y_in <= "10010001"; x_in <= "10010000"; z_correct<="0011000010010000";
        when 4369 => y_in <= "10010001"; x_in <= "10010001"; z_correct<="0011000000100001";
        when 4370 => y_in <= "10010001"; x_in <= "10010010"; z_correct<="0010111110110010";
        when 4371 => y_in <= "10010001"; x_in <= "10010011"; z_correct<="0010111101000011";
        when 4372 => y_in <= "10010001"; x_in <= "10010100"; z_correct<="0010111011010100";
        when 4373 => y_in <= "10010001"; x_in <= "10010101"; z_correct<="0010111001100101";
        when 4374 => y_in <= "10010001"; x_in <= "10010110"; z_correct<="0010110111110110";
        when 4375 => y_in <= "10010001"; x_in <= "10010111"; z_correct<="0010110110000111";
        when 4376 => y_in <= "10010001"; x_in <= "10011000"; z_correct<="0010110100011000";
        when 4377 => y_in <= "10010001"; x_in <= "10011001"; z_correct<="0010110010101001";
        when 4378 => y_in <= "10010001"; x_in <= "10011010"; z_correct<="0010110000111010";
        when 4379 => y_in <= "10010001"; x_in <= "10011011"; z_correct<="0010101111001011";
        when 4380 => y_in <= "10010001"; x_in <= "10011100"; z_correct<="0010101101011100";
        when 4381 => y_in <= "10010001"; x_in <= "10011101"; z_correct<="0010101011101101";
        when 4382 => y_in <= "10010001"; x_in <= "10011110"; z_correct<="0010101001111110";
        when 4383 => y_in <= "10010001"; x_in <= "10011111"; z_correct<="0010101000001111";
        when 4384 => y_in <= "10010001"; x_in <= "10100000"; z_correct<="0010100110100000";
        when 4385 => y_in <= "10010001"; x_in <= "10100001"; z_correct<="0010100100110001";
        when 4386 => y_in <= "10010001"; x_in <= "10100010"; z_correct<="0010100011000010";
        when 4387 => y_in <= "10010001"; x_in <= "10100011"; z_correct<="0010100001010011";
        when 4388 => y_in <= "10010001"; x_in <= "10100100"; z_correct<="0010011111100100";
        when 4389 => y_in <= "10010001"; x_in <= "10100101"; z_correct<="0010011101110101";
        when 4390 => y_in <= "10010001"; x_in <= "10100110"; z_correct<="0010011100000110";
        when 4391 => y_in <= "10010001"; x_in <= "10100111"; z_correct<="0010011010010111";
        when 4392 => y_in <= "10010001"; x_in <= "10101000"; z_correct<="0010011000101000";
        when 4393 => y_in <= "10010001"; x_in <= "10101001"; z_correct<="0010010110111001";
        when 4394 => y_in <= "10010001"; x_in <= "10101010"; z_correct<="0010010101001010";
        when 4395 => y_in <= "10010001"; x_in <= "10101011"; z_correct<="0010010011011011";
        when 4396 => y_in <= "10010001"; x_in <= "10101100"; z_correct<="0010010001101100";
        when 4397 => y_in <= "10010001"; x_in <= "10101101"; z_correct<="0010001111111101";
        when 4398 => y_in <= "10010001"; x_in <= "10101110"; z_correct<="0010001110001110";
        when 4399 => y_in <= "10010001"; x_in <= "10101111"; z_correct<="0010001100011111";
        when 4400 => y_in <= "10010001"; x_in <= "10110000"; z_correct<="0010001010110000";
        when 4401 => y_in <= "10010001"; x_in <= "10110001"; z_correct<="0010001001000001";
        when 4402 => y_in <= "10010001"; x_in <= "10110010"; z_correct<="0010000111010010";
        when 4403 => y_in <= "10010001"; x_in <= "10110011"; z_correct<="0010000101100011";
        when 4404 => y_in <= "10010001"; x_in <= "10110100"; z_correct<="0010000011110100";
        when 4405 => y_in <= "10010001"; x_in <= "10110101"; z_correct<="0010000010000101";
        when 4406 => y_in <= "10010001"; x_in <= "10110110"; z_correct<="0010000000010110";
        when 4407 => y_in <= "10010001"; x_in <= "10110111"; z_correct<="0001111110100111";
        when 4408 => y_in <= "10010001"; x_in <= "10111000"; z_correct<="0001111100111000";
        when 4409 => y_in <= "10010001"; x_in <= "10111001"; z_correct<="0001111011001001";
        when 4410 => y_in <= "10010001"; x_in <= "10111010"; z_correct<="0001111001011010";
        when 4411 => y_in <= "10010001"; x_in <= "10111011"; z_correct<="0001110111101011";
        when 4412 => y_in <= "10010001"; x_in <= "10111100"; z_correct<="0001110101111100";
        when 4413 => y_in <= "10010001"; x_in <= "10111101"; z_correct<="0001110100001101";
        when 4414 => y_in <= "10010001"; x_in <= "10111110"; z_correct<="0001110010011110";
        when 4415 => y_in <= "10010001"; x_in <= "10111111"; z_correct<="0001110000101111";
        when 4416 => y_in <= "10010001"; x_in <= "11000000"; z_correct<="0001101111000000";
        when 4417 => y_in <= "10010001"; x_in <= "11000001"; z_correct<="0001101101010001";
        when 4418 => y_in <= "10010001"; x_in <= "11000010"; z_correct<="0001101011100010";
        when 4419 => y_in <= "10010001"; x_in <= "11000011"; z_correct<="0001101001110011";
        when 4420 => y_in <= "10010001"; x_in <= "11000100"; z_correct<="0001101000000100";
        when 4421 => y_in <= "10010001"; x_in <= "11000101"; z_correct<="0001100110010101";
        when 4422 => y_in <= "10010001"; x_in <= "11000110"; z_correct<="0001100100100110";
        when 4423 => y_in <= "10010001"; x_in <= "11000111"; z_correct<="0001100010110111";
        when 4424 => y_in <= "10010001"; x_in <= "11001000"; z_correct<="0001100001001000";
        when 4425 => y_in <= "10010001"; x_in <= "11001001"; z_correct<="0001011111011001";
        when 4426 => y_in <= "10010001"; x_in <= "11001010"; z_correct<="0001011101101010";
        when 4427 => y_in <= "10010001"; x_in <= "11001011"; z_correct<="0001011011111011";
        when 4428 => y_in <= "10010001"; x_in <= "11001100"; z_correct<="0001011010001100";
        when 4429 => y_in <= "10010001"; x_in <= "11001101"; z_correct<="0001011000011101";
        when 4430 => y_in <= "10010001"; x_in <= "11001110"; z_correct<="0001010110101110";
        when 4431 => y_in <= "10010001"; x_in <= "11001111"; z_correct<="0001010100111111";
        when 4432 => y_in <= "10010001"; x_in <= "11010000"; z_correct<="0001010011010000";
        when 4433 => y_in <= "10010001"; x_in <= "11010001"; z_correct<="0001010001100001";
        when 4434 => y_in <= "10010001"; x_in <= "11010010"; z_correct<="0001001111110010";
        when 4435 => y_in <= "10010001"; x_in <= "11010011"; z_correct<="0001001110000011";
        when 4436 => y_in <= "10010001"; x_in <= "11010100"; z_correct<="0001001100010100";
        when 4437 => y_in <= "10010001"; x_in <= "11010101"; z_correct<="0001001010100101";
        when 4438 => y_in <= "10010001"; x_in <= "11010110"; z_correct<="0001001000110110";
        when 4439 => y_in <= "10010001"; x_in <= "11010111"; z_correct<="0001000111000111";
        when 4440 => y_in <= "10010001"; x_in <= "11011000"; z_correct<="0001000101011000";
        when 4441 => y_in <= "10010001"; x_in <= "11011001"; z_correct<="0001000011101001";
        when 4442 => y_in <= "10010001"; x_in <= "11011010"; z_correct<="0001000001111010";
        when 4443 => y_in <= "10010001"; x_in <= "11011011"; z_correct<="0001000000001011";
        when 4444 => y_in <= "10010001"; x_in <= "11011100"; z_correct<="0000111110011100";
        when 4445 => y_in <= "10010001"; x_in <= "11011101"; z_correct<="0000111100101101";
        when 4446 => y_in <= "10010001"; x_in <= "11011110"; z_correct<="0000111010111110";
        when 4447 => y_in <= "10010001"; x_in <= "11011111"; z_correct<="0000111001001111";
        when 4448 => y_in <= "10010001"; x_in <= "11100000"; z_correct<="0000110111100000";
        when 4449 => y_in <= "10010001"; x_in <= "11100001"; z_correct<="0000110101110001";
        when 4450 => y_in <= "10010001"; x_in <= "11100010"; z_correct<="0000110100000010";
        when 4451 => y_in <= "10010001"; x_in <= "11100011"; z_correct<="0000110010010011";
        when 4452 => y_in <= "10010001"; x_in <= "11100100"; z_correct<="0000110000100100";
        when 4453 => y_in <= "10010001"; x_in <= "11100101"; z_correct<="0000101110110101";
        when 4454 => y_in <= "10010001"; x_in <= "11100110"; z_correct<="0000101101000110";
        when 4455 => y_in <= "10010001"; x_in <= "11100111"; z_correct<="0000101011010111";
        when 4456 => y_in <= "10010001"; x_in <= "11101000"; z_correct<="0000101001101000";
        when 4457 => y_in <= "10010001"; x_in <= "11101001"; z_correct<="0000100111111001";
        when 4458 => y_in <= "10010001"; x_in <= "11101010"; z_correct<="0000100110001010";
        when 4459 => y_in <= "10010001"; x_in <= "11101011"; z_correct<="0000100100011011";
        when 4460 => y_in <= "10010001"; x_in <= "11101100"; z_correct<="0000100010101100";
        when 4461 => y_in <= "10010001"; x_in <= "11101101"; z_correct<="0000100000111101";
        when 4462 => y_in <= "10010001"; x_in <= "11101110"; z_correct<="0000011111001110";
        when 4463 => y_in <= "10010001"; x_in <= "11101111"; z_correct<="0000011101011111";
        when 4464 => y_in <= "10010001"; x_in <= "11110000"; z_correct<="0000011011110000";
        when 4465 => y_in <= "10010001"; x_in <= "11110001"; z_correct<="0000011010000001";
        when 4466 => y_in <= "10010001"; x_in <= "11110010"; z_correct<="0000011000010010";
        when 4467 => y_in <= "10010001"; x_in <= "11110011"; z_correct<="0000010110100011";
        when 4468 => y_in <= "10010001"; x_in <= "11110100"; z_correct<="0000010100110100";
        when 4469 => y_in <= "10010001"; x_in <= "11110101"; z_correct<="0000010011000101";
        when 4470 => y_in <= "10010001"; x_in <= "11110110"; z_correct<="0000010001010110";
        when 4471 => y_in <= "10010001"; x_in <= "11110111"; z_correct<="0000001111100111";
        when 4472 => y_in <= "10010001"; x_in <= "11111000"; z_correct<="0000001101111000";
        when 4473 => y_in <= "10010001"; x_in <= "11111001"; z_correct<="0000001100001001";
        when 4474 => y_in <= "10010001"; x_in <= "11111010"; z_correct<="0000001010011010";
        when 4475 => y_in <= "10010001"; x_in <= "11111011"; z_correct<="0000001000101011";
        when 4476 => y_in <= "10010001"; x_in <= "11111100"; z_correct<="0000000110111100";
        when 4477 => y_in <= "10010001"; x_in <= "11111101"; z_correct<="0000000101001101";
        when 4478 => y_in <= "10010001"; x_in <= "11111110"; z_correct<="0000000011011110";
        when 4479 => y_in <= "10010001"; x_in <= "11111111"; z_correct<="0000000001101111";
        when 4480 => y_in <= "10010001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 4481 => y_in <= "10010001"; x_in <= "00000001"; z_correct<="1111111110010001";
        when 4482 => y_in <= "10010001"; x_in <= "00000010"; z_correct<="1111111100100010";
        when 4483 => y_in <= "10010001"; x_in <= "00000011"; z_correct<="1111111010110011";
        when 4484 => y_in <= "10010001"; x_in <= "00000100"; z_correct<="1111111001000100";
        when 4485 => y_in <= "10010001"; x_in <= "00000101"; z_correct<="1111110111010101";
        when 4486 => y_in <= "10010001"; x_in <= "00000110"; z_correct<="1111110101100110";
        when 4487 => y_in <= "10010001"; x_in <= "00000111"; z_correct<="1111110011110111";
        when 4488 => y_in <= "10010001"; x_in <= "00001000"; z_correct<="1111110010001000";
        when 4489 => y_in <= "10010001"; x_in <= "00001001"; z_correct<="1111110000011001";
        when 4490 => y_in <= "10010001"; x_in <= "00001010"; z_correct<="1111101110101010";
        when 4491 => y_in <= "10010001"; x_in <= "00001011"; z_correct<="1111101100111011";
        when 4492 => y_in <= "10010001"; x_in <= "00001100"; z_correct<="1111101011001100";
        when 4493 => y_in <= "10010001"; x_in <= "00001101"; z_correct<="1111101001011101";
        when 4494 => y_in <= "10010001"; x_in <= "00001110"; z_correct<="1111100111101110";
        when 4495 => y_in <= "10010001"; x_in <= "00001111"; z_correct<="1111100101111111";
        when 4496 => y_in <= "10010001"; x_in <= "00010000"; z_correct<="1111100100010000";
        when 4497 => y_in <= "10010001"; x_in <= "00010001"; z_correct<="1111100010100001";
        when 4498 => y_in <= "10010001"; x_in <= "00010010"; z_correct<="1111100000110010";
        when 4499 => y_in <= "10010001"; x_in <= "00010011"; z_correct<="1111011111000011";
        when 4500 => y_in <= "10010001"; x_in <= "00010100"; z_correct<="1111011101010100";
        when 4501 => y_in <= "10010001"; x_in <= "00010101"; z_correct<="1111011011100101";
        when 4502 => y_in <= "10010001"; x_in <= "00010110"; z_correct<="1111011001110110";
        when 4503 => y_in <= "10010001"; x_in <= "00010111"; z_correct<="1111011000000111";
        when 4504 => y_in <= "10010001"; x_in <= "00011000"; z_correct<="1111010110011000";
        when 4505 => y_in <= "10010001"; x_in <= "00011001"; z_correct<="1111010100101001";
        when 4506 => y_in <= "10010001"; x_in <= "00011010"; z_correct<="1111010010111010";
        when 4507 => y_in <= "10010001"; x_in <= "00011011"; z_correct<="1111010001001011";
        when 4508 => y_in <= "10010001"; x_in <= "00011100"; z_correct<="1111001111011100";
        when 4509 => y_in <= "10010001"; x_in <= "00011101"; z_correct<="1111001101101101";
        when 4510 => y_in <= "10010001"; x_in <= "00011110"; z_correct<="1111001011111110";
        when 4511 => y_in <= "10010001"; x_in <= "00011111"; z_correct<="1111001010001111";
        when 4512 => y_in <= "10010001"; x_in <= "00100000"; z_correct<="1111001000100000";
        when 4513 => y_in <= "10010001"; x_in <= "00100001"; z_correct<="1111000110110001";
        when 4514 => y_in <= "10010001"; x_in <= "00100010"; z_correct<="1111000101000010";
        when 4515 => y_in <= "10010001"; x_in <= "00100011"; z_correct<="1111000011010011";
        when 4516 => y_in <= "10010001"; x_in <= "00100100"; z_correct<="1111000001100100";
        when 4517 => y_in <= "10010001"; x_in <= "00100101"; z_correct<="1110111111110101";
        when 4518 => y_in <= "10010001"; x_in <= "00100110"; z_correct<="1110111110000110";
        when 4519 => y_in <= "10010001"; x_in <= "00100111"; z_correct<="1110111100010111";
        when 4520 => y_in <= "10010001"; x_in <= "00101000"; z_correct<="1110111010101000";
        when 4521 => y_in <= "10010001"; x_in <= "00101001"; z_correct<="1110111000111001";
        when 4522 => y_in <= "10010001"; x_in <= "00101010"; z_correct<="1110110111001010";
        when 4523 => y_in <= "10010001"; x_in <= "00101011"; z_correct<="1110110101011011";
        when 4524 => y_in <= "10010001"; x_in <= "00101100"; z_correct<="1110110011101100";
        when 4525 => y_in <= "10010001"; x_in <= "00101101"; z_correct<="1110110001111101";
        when 4526 => y_in <= "10010001"; x_in <= "00101110"; z_correct<="1110110000001110";
        when 4527 => y_in <= "10010001"; x_in <= "00101111"; z_correct<="1110101110011111";
        when 4528 => y_in <= "10010001"; x_in <= "00110000"; z_correct<="1110101100110000";
        when 4529 => y_in <= "10010001"; x_in <= "00110001"; z_correct<="1110101011000001";
        when 4530 => y_in <= "10010001"; x_in <= "00110010"; z_correct<="1110101001010010";
        when 4531 => y_in <= "10010001"; x_in <= "00110011"; z_correct<="1110100111100011";
        when 4532 => y_in <= "10010001"; x_in <= "00110100"; z_correct<="1110100101110100";
        when 4533 => y_in <= "10010001"; x_in <= "00110101"; z_correct<="1110100100000101";
        when 4534 => y_in <= "10010001"; x_in <= "00110110"; z_correct<="1110100010010110";
        when 4535 => y_in <= "10010001"; x_in <= "00110111"; z_correct<="1110100000100111";
        when 4536 => y_in <= "10010001"; x_in <= "00111000"; z_correct<="1110011110111000";
        when 4537 => y_in <= "10010001"; x_in <= "00111001"; z_correct<="1110011101001001";
        when 4538 => y_in <= "10010001"; x_in <= "00111010"; z_correct<="1110011011011010";
        when 4539 => y_in <= "10010001"; x_in <= "00111011"; z_correct<="1110011001101011";
        when 4540 => y_in <= "10010001"; x_in <= "00111100"; z_correct<="1110010111111100";
        when 4541 => y_in <= "10010001"; x_in <= "00111101"; z_correct<="1110010110001101";
        when 4542 => y_in <= "10010001"; x_in <= "00111110"; z_correct<="1110010100011110";
        when 4543 => y_in <= "10010001"; x_in <= "00111111"; z_correct<="1110010010101111";
        when 4544 => y_in <= "10010001"; x_in <= "01000000"; z_correct<="1110010001000000";
        when 4545 => y_in <= "10010001"; x_in <= "01000001"; z_correct<="1110001111010001";
        when 4546 => y_in <= "10010001"; x_in <= "01000010"; z_correct<="1110001101100010";
        when 4547 => y_in <= "10010001"; x_in <= "01000011"; z_correct<="1110001011110011";
        when 4548 => y_in <= "10010001"; x_in <= "01000100"; z_correct<="1110001010000100";
        when 4549 => y_in <= "10010001"; x_in <= "01000101"; z_correct<="1110001000010101";
        when 4550 => y_in <= "10010001"; x_in <= "01000110"; z_correct<="1110000110100110";
        when 4551 => y_in <= "10010001"; x_in <= "01000111"; z_correct<="1110000100110111";
        when 4552 => y_in <= "10010001"; x_in <= "01001000"; z_correct<="1110000011001000";
        when 4553 => y_in <= "10010001"; x_in <= "01001001"; z_correct<="1110000001011001";
        when 4554 => y_in <= "10010001"; x_in <= "01001010"; z_correct<="1101111111101010";
        when 4555 => y_in <= "10010001"; x_in <= "01001011"; z_correct<="1101111101111011";
        when 4556 => y_in <= "10010001"; x_in <= "01001100"; z_correct<="1101111100001100";
        when 4557 => y_in <= "10010001"; x_in <= "01001101"; z_correct<="1101111010011101";
        when 4558 => y_in <= "10010001"; x_in <= "01001110"; z_correct<="1101111000101110";
        when 4559 => y_in <= "10010001"; x_in <= "01001111"; z_correct<="1101110110111111";
        when 4560 => y_in <= "10010001"; x_in <= "01010000"; z_correct<="1101110101010000";
        when 4561 => y_in <= "10010001"; x_in <= "01010001"; z_correct<="1101110011100001";
        when 4562 => y_in <= "10010001"; x_in <= "01010010"; z_correct<="1101110001110010";
        when 4563 => y_in <= "10010001"; x_in <= "01010011"; z_correct<="1101110000000011";
        when 4564 => y_in <= "10010001"; x_in <= "01010100"; z_correct<="1101101110010100";
        when 4565 => y_in <= "10010001"; x_in <= "01010101"; z_correct<="1101101100100101";
        when 4566 => y_in <= "10010001"; x_in <= "01010110"; z_correct<="1101101010110110";
        when 4567 => y_in <= "10010001"; x_in <= "01010111"; z_correct<="1101101001000111";
        when 4568 => y_in <= "10010001"; x_in <= "01011000"; z_correct<="1101100111011000";
        when 4569 => y_in <= "10010001"; x_in <= "01011001"; z_correct<="1101100101101001";
        when 4570 => y_in <= "10010001"; x_in <= "01011010"; z_correct<="1101100011111010";
        when 4571 => y_in <= "10010001"; x_in <= "01011011"; z_correct<="1101100010001011";
        when 4572 => y_in <= "10010001"; x_in <= "01011100"; z_correct<="1101100000011100";
        when 4573 => y_in <= "10010001"; x_in <= "01011101"; z_correct<="1101011110101101";
        when 4574 => y_in <= "10010001"; x_in <= "01011110"; z_correct<="1101011100111110";
        when 4575 => y_in <= "10010001"; x_in <= "01011111"; z_correct<="1101011011001111";
        when 4576 => y_in <= "10010001"; x_in <= "01100000"; z_correct<="1101011001100000";
        when 4577 => y_in <= "10010001"; x_in <= "01100001"; z_correct<="1101010111110001";
        when 4578 => y_in <= "10010001"; x_in <= "01100010"; z_correct<="1101010110000010";
        when 4579 => y_in <= "10010001"; x_in <= "01100011"; z_correct<="1101010100010011";
        when 4580 => y_in <= "10010001"; x_in <= "01100100"; z_correct<="1101010010100100";
        when 4581 => y_in <= "10010001"; x_in <= "01100101"; z_correct<="1101010000110101";
        when 4582 => y_in <= "10010001"; x_in <= "01100110"; z_correct<="1101001111000110";
        when 4583 => y_in <= "10010001"; x_in <= "01100111"; z_correct<="1101001101010111";
        when 4584 => y_in <= "10010001"; x_in <= "01101000"; z_correct<="1101001011101000";
        when 4585 => y_in <= "10010001"; x_in <= "01101001"; z_correct<="1101001001111001";
        when 4586 => y_in <= "10010001"; x_in <= "01101010"; z_correct<="1101001000001010";
        when 4587 => y_in <= "10010001"; x_in <= "01101011"; z_correct<="1101000110011011";
        when 4588 => y_in <= "10010001"; x_in <= "01101100"; z_correct<="1101000100101100";
        when 4589 => y_in <= "10010001"; x_in <= "01101101"; z_correct<="1101000010111101";
        when 4590 => y_in <= "10010001"; x_in <= "01101110"; z_correct<="1101000001001110";
        when 4591 => y_in <= "10010001"; x_in <= "01101111"; z_correct<="1100111111011111";
        when 4592 => y_in <= "10010001"; x_in <= "01110000"; z_correct<="1100111101110000";
        when 4593 => y_in <= "10010001"; x_in <= "01110001"; z_correct<="1100111100000001";
        when 4594 => y_in <= "10010001"; x_in <= "01110010"; z_correct<="1100111010010010";
        when 4595 => y_in <= "10010001"; x_in <= "01110011"; z_correct<="1100111000100011";
        when 4596 => y_in <= "10010001"; x_in <= "01110100"; z_correct<="1100110110110100";
        when 4597 => y_in <= "10010001"; x_in <= "01110101"; z_correct<="1100110101000101";
        when 4598 => y_in <= "10010001"; x_in <= "01110110"; z_correct<="1100110011010110";
        when 4599 => y_in <= "10010001"; x_in <= "01110111"; z_correct<="1100110001100111";
        when 4600 => y_in <= "10010001"; x_in <= "01111000"; z_correct<="1100101111111000";
        when 4601 => y_in <= "10010001"; x_in <= "01111001"; z_correct<="1100101110001001";
        when 4602 => y_in <= "10010001"; x_in <= "01111010"; z_correct<="1100101100011010";
        when 4603 => y_in <= "10010001"; x_in <= "01111011"; z_correct<="1100101010101011";
        when 4604 => y_in <= "10010001"; x_in <= "01111100"; z_correct<="1100101000111100";
        when 4605 => y_in <= "10010001"; x_in <= "01111101"; z_correct<="1100100111001101";
        when 4606 => y_in <= "10010001"; x_in <= "01111110"; z_correct<="1100100101011110";
        when 4607 => y_in <= "10010001"; x_in <= "01111111"; z_correct<="1100100011101111";
        when 4608 => y_in <= "10010010"; x_in <= "10000000"; z_correct<="0011011100000000";
        when 4609 => y_in <= "10010010"; x_in <= "10000001"; z_correct<="0011011010010010";
        when 4610 => y_in <= "10010010"; x_in <= "10000010"; z_correct<="0011011000100100";
        when 4611 => y_in <= "10010010"; x_in <= "10000011"; z_correct<="0011010110110110";
        when 4612 => y_in <= "10010010"; x_in <= "10000100"; z_correct<="0011010101001000";
        when 4613 => y_in <= "10010010"; x_in <= "10000101"; z_correct<="0011010011011010";
        when 4614 => y_in <= "10010010"; x_in <= "10000110"; z_correct<="0011010001101100";
        when 4615 => y_in <= "10010010"; x_in <= "10000111"; z_correct<="0011001111111110";
        when 4616 => y_in <= "10010010"; x_in <= "10001000"; z_correct<="0011001110010000";
        when 4617 => y_in <= "10010010"; x_in <= "10001001"; z_correct<="0011001100100010";
        when 4618 => y_in <= "10010010"; x_in <= "10001010"; z_correct<="0011001010110100";
        when 4619 => y_in <= "10010010"; x_in <= "10001011"; z_correct<="0011001001000110";
        when 4620 => y_in <= "10010010"; x_in <= "10001100"; z_correct<="0011000111011000";
        when 4621 => y_in <= "10010010"; x_in <= "10001101"; z_correct<="0011000101101010";
        when 4622 => y_in <= "10010010"; x_in <= "10001110"; z_correct<="0011000011111100";
        when 4623 => y_in <= "10010010"; x_in <= "10001111"; z_correct<="0011000010001110";
        when 4624 => y_in <= "10010010"; x_in <= "10010000"; z_correct<="0011000000100000";
        when 4625 => y_in <= "10010010"; x_in <= "10010001"; z_correct<="0010111110110010";
        when 4626 => y_in <= "10010010"; x_in <= "10010010"; z_correct<="0010111101000100";
        when 4627 => y_in <= "10010010"; x_in <= "10010011"; z_correct<="0010111011010110";
        when 4628 => y_in <= "10010010"; x_in <= "10010100"; z_correct<="0010111001101000";
        when 4629 => y_in <= "10010010"; x_in <= "10010101"; z_correct<="0010110111111010";
        when 4630 => y_in <= "10010010"; x_in <= "10010110"; z_correct<="0010110110001100";
        when 4631 => y_in <= "10010010"; x_in <= "10010111"; z_correct<="0010110100011110";
        when 4632 => y_in <= "10010010"; x_in <= "10011000"; z_correct<="0010110010110000";
        when 4633 => y_in <= "10010010"; x_in <= "10011001"; z_correct<="0010110001000010";
        when 4634 => y_in <= "10010010"; x_in <= "10011010"; z_correct<="0010101111010100";
        when 4635 => y_in <= "10010010"; x_in <= "10011011"; z_correct<="0010101101100110";
        when 4636 => y_in <= "10010010"; x_in <= "10011100"; z_correct<="0010101011111000";
        when 4637 => y_in <= "10010010"; x_in <= "10011101"; z_correct<="0010101010001010";
        when 4638 => y_in <= "10010010"; x_in <= "10011110"; z_correct<="0010101000011100";
        when 4639 => y_in <= "10010010"; x_in <= "10011111"; z_correct<="0010100110101110";
        when 4640 => y_in <= "10010010"; x_in <= "10100000"; z_correct<="0010100101000000";
        when 4641 => y_in <= "10010010"; x_in <= "10100001"; z_correct<="0010100011010010";
        when 4642 => y_in <= "10010010"; x_in <= "10100010"; z_correct<="0010100001100100";
        when 4643 => y_in <= "10010010"; x_in <= "10100011"; z_correct<="0010011111110110";
        when 4644 => y_in <= "10010010"; x_in <= "10100100"; z_correct<="0010011110001000";
        when 4645 => y_in <= "10010010"; x_in <= "10100101"; z_correct<="0010011100011010";
        when 4646 => y_in <= "10010010"; x_in <= "10100110"; z_correct<="0010011010101100";
        when 4647 => y_in <= "10010010"; x_in <= "10100111"; z_correct<="0010011000111110";
        when 4648 => y_in <= "10010010"; x_in <= "10101000"; z_correct<="0010010111010000";
        when 4649 => y_in <= "10010010"; x_in <= "10101001"; z_correct<="0010010101100010";
        when 4650 => y_in <= "10010010"; x_in <= "10101010"; z_correct<="0010010011110100";
        when 4651 => y_in <= "10010010"; x_in <= "10101011"; z_correct<="0010010010000110";
        when 4652 => y_in <= "10010010"; x_in <= "10101100"; z_correct<="0010010000011000";
        when 4653 => y_in <= "10010010"; x_in <= "10101101"; z_correct<="0010001110101010";
        when 4654 => y_in <= "10010010"; x_in <= "10101110"; z_correct<="0010001100111100";
        when 4655 => y_in <= "10010010"; x_in <= "10101111"; z_correct<="0010001011001110";
        when 4656 => y_in <= "10010010"; x_in <= "10110000"; z_correct<="0010001001100000";
        when 4657 => y_in <= "10010010"; x_in <= "10110001"; z_correct<="0010000111110010";
        when 4658 => y_in <= "10010010"; x_in <= "10110010"; z_correct<="0010000110000100";
        when 4659 => y_in <= "10010010"; x_in <= "10110011"; z_correct<="0010000100010110";
        when 4660 => y_in <= "10010010"; x_in <= "10110100"; z_correct<="0010000010101000";
        when 4661 => y_in <= "10010010"; x_in <= "10110101"; z_correct<="0010000000111010";
        when 4662 => y_in <= "10010010"; x_in <= "10110110"; z_correct<="0001111111001100";
        when 4663 => y_in <= "10010010"; x_in <= "10110111"; z_correct<="0001111101011110";
        when 4664 => y_in <= "10010010"; x_in <= "10111000"; z_correct<="0001111011110000";
        when 4665 => y_in <= "10010010"; x_in <= "10111001"; z_correct<="0001111010000010";
        when 4666 => y_in <= "10010010"; x_in <= "10111010"; z_correct<="0001111000010100";
        when 4667 => y_in <= "10010010"; x_in <= "10111011"; z_correct<="0001110110100110";
        when 4668 => y_in <= "10010010"; x_in <= "10111100"; z_correct<="0001110100111000";
        when 4669 => y_in <= "10010010"; x_in <= "10111101"; z_correct<="0001110011001010";
        when 4670 => y_in <= "10010010"; x_in <= "10111110"; z_correct<="0001110001011100";
        when 4671 => y_in <= "10010010"; x_in <= "10111111"; z_correct<="0001101111101110";
        when 4672 => y_in <= "10010010"; x_in <= "11000000"; z_correct<="0001101110000000";
        when 4673 => y_in <= "10010010"; x_in <= "11000001"; z_correct<="0001101100010010";
        when 4674 => y_in <= "10010010"; x_in <= "11000010"; z_correct<="0001101010100100";
        when 4675 => y_in <= "10010010"; x_in <= "11000011"; z_correct<="0001101000110110";
        when 4676 => y_in <= "10010010"; x_in <= "11000100"; z_correct<="0001100111001000";
        when 4677 => y_in <= "10010010"; x_in <= "11000101"; z_correct<="0001100101011010";
        when 4678 => y_in <= "10010010"; x_in <= "11000110"; z_correct<="0001100011101100";
        when 4679 => y_in <= "10010010"; x_in <= "11000111"; z_correct<="0001100001111110";
        when 4680 => y_in <= "10010010"; x_in <= "11001000"; z_correct<="0001100000010000";
        when 4681 => y_in <= "10010010"; x_in <= "11001001"; z_correct<="0001011110100010";
        when 4682 => y_in <= "10010010"; x_in <= "11001010"; z_correct<="0001011100110100";
        when 4683 => y_in <= "10010010"; x_in <= "11001011"; z_correct<="0001011011000110";
        when 4684 => y_in <= "10010010"; x_in <= "11001100"; z_correct<="0001011001011000";
        when 4685 => y_in <= "10010010"; x_in <= "11001101"; z_correct<="0001010111101010";
        when 4686 => y_in <= "10010010"; x_in <= "11001110"; z_correct<="0001010101111100";
        when 4687 => y_in <= "10010010"; x_in <= "11001111"; z_correct<="0001010100001110";
        when 4688 => y_in <= "10010010"; x_in <= "11010000"; z_correct<="0001010010100000";
        when 4689 => y_in <= "10010010"; x_in <= "11010001"; z_correct<="0001010000110010";
        when 4690 => y_in <= "10010010"; x_in <= "11010010"; z_correct<="0001001111000100";
        when 4691 => y_in <= "10010010"; x_in <= "11010011"; z_correct<="0001001101010110";
        when 4692 => y_in <= "10010010"; x_in <= "11010100"; z_correct<="0001001011101000";
        when 4693 => y_in <= "10010010"; x_in <= "11010101"; z_correct<="0001001001111010";
        when 4694 => y_in <= "10010010"; x_in <= "11010110"; z_correct<="0001001000001100";
        when 4695 => y_in <= "10010010"; x_in <= "11010111"; z_correct<="0001000110011110";
        when 4696 => y_in <= "10010010"; x_in <= "11011000"; z_correct<="0001000100110000";
        when 4697 => y_in <= "10010010"; x_in <= "11011001"; z_correct<="0001000011000010";
        when 4698 => y_in <= "10010010"; x_in <= "11011010"; z_correct<="0001000001010100";
        when 4699 => y_in <= "10010010"; x_in <= "11011011"; z_correct<="0000111111100110";
        when 4700 => y_in <= "10010010"; x_in <= "11011100"; z_correct<="0000111101111000";
        when 4701 => y_in <= "10010010"; x_in <= "11011101"; z_correct<="0000111100001010";
        when 4702 => y_in <= "10010010"; x_in <= "11011110"; z_correct<="0000111010011100";
        when 4703 => y_in <= "10010010"; x_in <= "11011111"; z_correct<="0000111000101110";
        when 4704 => y_in <= "10010010"; x_in <= "11100000"; z_correct<="0000110111000000";
        when 4705 => y_in <= "10010010"; x_in <= "11100001"; z_correct<="0000110101010010";
        when 4706 => y_in <= "10010010"; x_in <= "11100010"; z_correct<="0000110011100100";
        when 4707 => y_in <= "10010010"; x_in <= "11100011"; z_correct<="0000110001110110";
        when 4708 => y_in <= "10010010"; x_in <= "11100100"; z_correct<="0000110000001000";
        when 4709 => y_in <= "10010010"; x_in <= "11100101"; z_correct<="0000101110011010";
        when 4710 => y_in <= "10010010"; x_in <= "11100110"; z_correct<="0000101100101100";
        when 4711 => y_in <= "10010010"; x_in <= "11100111"; z_correct<="0000101010111110";
        when 4712 => y_in <= "10010010"; x_in <= "11101000"; z_correct<="0000101001010000";
        when 4713 => y_in <= "10010010"; x_in <= "11101001"; z_correct<="0000100111100010";
        when 4714 => y_in <= "10010010"; x_in <= "11101010"; z_correct<="0000100101110100";
        when 4715 => y_in <= "10010010"; x_in <= "11101011"; z_correct<="0000100100000110";
        when 4716 => y_in <= "10010010"; x_in <= "11101100"; z_correct<="0000100010011000";
        when 4717 => y_in <= "10010010"; x_in <= "11101101"; z_correct<="0000100000101010";
        when 4718 => y_in <= "10010010"; x_in <= "11101110"; z_correct<="0000011110111100";
        when 4719 => y_in <= "10010010"; x_in <= "11101111"; z_correct<="0000011101001110";
        when 4720 => y_in <= "10010010"; x_in <= "11110000"; z_correct<="0000011011100000";
        when 4721 => y_in <= "10010010"; x_in <= "11110001"; z_correct<="0000011001110010";
        when 4722 => y_in <= "10010010"; x_in <= "11110010"; z_correct<="0000011000000100";
        when 4723 => y_in <= "10010010"; x_in <= "11110011"; z_correct<="0000010110010110";
        when 4724 => y_in <= "10010010"; x_in <= "11110100"; z_correct<="0000010100101000";
        when 4725 => y_in <= "10010010"; x_in <= "11110101"; z_correct<="0000010010111010";
        when 4726 => y_in <= "10010010"; x_in <= "11110110"; z_correct<="0000010001001100";
        when 4727 => y_in <= "10010010"; x_in <= "11110111"; z_correct<="0000001111011110";
        when 4728 => y_in <= "10010010"; x_in <= "11111000"; z_correct<="0000001101110000";
        when 4729 => y_in <= "10010010"; x_in <= "11111001"; z_correct<="0000001100000010";
        when 4730 => y_in <= "10010010"; x_in <= "11111010"; z_correct<="0000001010010100";
        when 4731 => y_in <= "10010010"; x_in <= "11111011"; z_correct<="0000001000100110";
        when 4732 => y_in <= "10010010"; x_in <= "11111100"; z_correct<="0000000110111000";
        when 4733 => y_in <= "10010010"; x_in <= "11111101"; z_correct<="0000000101001010";
        when 4734 => y_in <= "10010010"; x_in <= "11111110"; z_correct<="0000000011011100";
        when 4735 => y_in <= "10010010"; x_in <= "11111111"; z_correct<="0000000001101110";
        when 4736 => y_in <= "10010010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 4737 => y_in <= "10010010"; x_in <= "00000001"; z_correct<="1111111110010010";
        when 4738 => y_in <= "10010010"; x_in <= "00000010"; z_correct<="1111111100100100";
        when 4739 => y_in <= "10010010"; x_in <= "00000011"; z_correct<="1111111010110110";
        when 4740 => y_in <= "10010010"; x_in <= "00000100"; z_correct<="1111111001001000";
        when 4741 => y_in <= "10010010"; x_in <= "00000101"; z_correct<="1111110111011010";
        when 4742 => y_in <= "10010010"; x_in <= "00000110"; z_correct<="1111110101101100";
        when 4743 => y_in <= "10010010"; x_in <= "00000111"; z_correct<="1111110011111110";
        when 4744 => y_in <= "10010010"; x_in <= "00001000"; z_correct<="1111110010010000";
        when 4745 => y_in <= "10010010"; x_in <= "00001001"; z_correct<="1111110000100010";
        when 4746 => y_in <= "10010010"; x_in <= "00001010"; z_correct<="1111101110110100";
        when 4747 => y_in <= "10010010"; x_in <= "00001011"; z_correct<="1111101101000110";
        when 4748 => y_in <= "10010010"; x_in <= "00001100"; z_correct<="1111101011011000";
        when 4749 => y_in <= "10010010"; x_in <= "00001101"; z_correct<="1111101001101010";
        when 4750 => y_in <= "10010010"; x_in <= "00001110"; z_correct<="1111100111111100";
        when 4751 => y_in <= "10010010"; x_in <= "00001111"; z_correct<="1111100110001110";
        when 4752 => y_in <= "10010010"; x_in <= "00010000"; z_correct<="1111100100100000";
        when 4753 => y_in <= "10010010"; x_in <= "00010001"; z_correct<="1111100010110010";
        when 4754 => y_in <= "10010010"; x_in <= "00010010"; z_correct<="1111100001000100";
        when 4755 => y_in <= "10010010"; x_in <= "00010011"; z_correct<="1111011111010110";
        when 4756 => y_in <= "10010010"; x_in <= "00010100"; z_correct<="1111011101101000";
        when 4757 => y_in <= "10010010"; x_in <= "00010101"; z_correct<="1111011011111010";
        when 4758 => y_in <= "10010010"; x_in <= "00010110"; z_correct<="1111011010001100";
        when 4759 => y_in <= "10010010"; x_in <= "00010111"; z_correct<="1111011000011110";
        when 4760 => y_in <= "10010010"; x_in <= "00011000"; z_correct<="1111010110110000";
        when 4761 => y_in <= "10010010"; x_in <= "00011001"; z_correct<="1111010101000010";
        when 4762 => y_in <= "10010010"; x_in <= "00011010"; z_correct<="1111010011010100";
        when 4763 => y_in <= "10010010"; x_in <= "00011011"; z_correct<="1111010001100110";
        when 4764 => y_in <= "10010010"; x_in <= "00011100"; z_correct<="1111001111111000";
        when 4765 => y_in <= "10010010"; x_in <= "00011101"; z_correct<="1111001110001010";
        when 4766 => y_in <= "10010010"; x_in <= "00011110"; z_correct<="1111001100011100";
        when 4767 => y_in <= "10010010"; x_in <= "00011111"; z_correct<="1111001010101110";
        when 4768 => y_in <= "10010010"; x_in <= "00100000"; z_correct<="1111001001000000";
        when 4769 => y_in <= "10010010"; x_in <= "00100001"; z_correct<="1111000111010010";
        when 4770 => y_in <= "10010010"; x_in <= "00100010"; z_correct<="1111000101100100";
        when 4771 => y_in <= "10010010"; x_in <= "00100011"; z_correct<="1111000011110110";
        when 4772 => y_in <= "10010010"; x_in <= "00100100"; z_correct<="1111000010001000";
        when 4773 => y_in <= "10010010"; x_in <= "00100101"; z_correct<="1111000000011010";
        when 4774 => y_in <= "10010010"; x_in <= "00100110"; z_correct<="1110111110101100";
        when 4775 => y_in <= "10010010"; x_in <= "00100111"; z_correct<="1110111100111110";
        when 4776 => y_in <= "10010010"; x_in <= "00101000"; z_correct<="1110111011010000";
        when 4777 => y_in <= "10010010"; x_in <= "00101001"; z_correct<="1110111001100010";
        when 4778 => y_in <= "10010010"; x_in <= "00101010"; z_correct<="1110110111110100";
        when 4779 => y_in <= "10010010"; x_in <= "00101011"; z_correct<="1110110110000110";
        when 4780 => y_in <= "10010010"; x_in <= "00101100"; z_correct<="1110110100011000";
        when 4781 => y_in <= "10010010"; x_in <= "00101101"; z_correct<="1110110010101010";
        when 4782 => y_in <= "10010010"; x_in <= "00101110"; z_correct<="1110110000111100";
        when 4783 => y_in <= "10010010"; x_in <= "00101111"; z_correct<="1110101111001110";
        when 4784 => y_in <= "10010010"; x_in <= "00110000"; z_correct<="1110101101100000";
        when 4785 => y_in <= "10010010"; x_in <= "00110001"; z_correct<="1110101011110010";
        when 4786 => y_in <= "10010010"; x_in <= "00110010"; z_correct<="1110101010000100";
        when 4787 => y_in <= "10010010"; x_in <= "00110011"; z_correct<="1110101000010110";
        when 4788 => y_in <= "10010010"; x_in <= "00110100"; z_correct<="1110100110101000";
        when 4789 => y_in <= "10010010"; x_in <= "00110101"; z_correct<="1110100100111010";
        when 4790 => y_in <= "10010010"; x_in <= "00110110"; z_correct<="1110100011001100";
        when 4791 => y_in <= "10010010"; x_in <= "00110111"; z_correct<="1110100001011110";
        when 4792 => y_in <= "10010010"; x_in <= "00111000"; z_correct<="1110011111110000";
        when 4793 => y_in <= "10010010"; x_in <= "00111001"; z_correct<="1110011110000010";
        when 4794 => y_in <= "10010010"; x_in <= "00111010"; z_correct<="1110011100010100";
        when 4795 => y_in <= "10010010"; x_in <= "00111011"; z_correct<="1110011010100110";
        when 4796 => y_in <= "10010010"; x_in <= "00111100"; z_correct<="1110011000111000";
        when 4797 => y_in <= "10010010"; x_in <= "00111101"; z_correct<="1110010111001010";
        when 4798 => y_in <= "10010010"; x_in <= "00111110"; z_correct<="1110010101011100";
        when 4799 => y_in <= "10010010"; x_in <= "00111111"; z_correct<="1110010011101110";
        when 4800 => y_in <= "10010010"; x_in <= "01000000"; z_correct<="1110010010000000";
        when 4801 => y_in <= "10010010"; x_in <= "01000001"; z_correct<="1110010000010010";
        when 4802 => y_in <= "10010010"; x_in <= "01000010"; z_correct<="1110001110100100";
        when 4803 => y_in <= "10010010"; x_in <= "01000011"; z_correct<="1110001100110110";
        when 4804 => y_in <= "10010010"; x_in <= "01000100"; z_correct<="1110001011001000";
        when 4805 => y_in <= "10010010"; x_in <= "01000101"; z_correct<="1110001001011010";
        when 4806 => y_in <= "10010010"; x_in <= "01000110"; z_correct<="1110000111101100";
        when 4807 => y_in <= "10010010"; x_in <= "01000111"; z_correct<="1110000101111110";
        when 4808 => y_in <= "10010010"; x_in <= "01001000"; z_correct<="1110000100010000";
        when 4809 => y_in <= "10010010"; x_in <= "01001001"; z_correct<="1110000010100010";
        when 4810 => y_in <= "10010010"; x_in <= "01001010"; z_correct<="1110000000110100";
        when 4811 => y_in <= "10010010"; x_in <= "01001011"; z_correct<="1101111111000110";
        when 4812 => y_in <= "10010010"; x_in <= "01001100"; z_correct<="1101111101011000";
        when 4813 => y_in <= "10010010"; x_in <= "01001101"; z_correct<="1101111011101010";
        when 4814 => y_in <= "10010010"; x_in <= "01001110"; z_correct<="1101111001111100";
        when 4815 => y_in <= "10010010"; x_in <= "01001111"; z_correct<="1101111000001110";
        when 4816 => y_in <= "10010010"; x_in <= "01010000"; z_correct<="1101110110100000";
        when 4817 => y_in <= "10010010"; x_in <= "01010001"; z_correct<="1101110100110010";
        when 4818 => y_in <= "10010010"; x_in <= "01010010"; z_correct<="1101110011000100";
        when 4819 => y_in <= "10010010"; x_in <= "01010011"; z_correct<="1101110001010110";
        when 4820 => y_in <= "10010010"; x_in <= "01010100"; z_correct<="1101101111101000";
        when 4821 => y_in <= "10010010"; x_in <= "01010101"; z_correct<="1101101101111010";
        when 4822 => y_in <= "10010010"; x_in <= "01010110"; z_correct<="1101101100001100";
        when 4823 => y_in <= "10010010"; x_in <= "01010111"; z_correct<="1101101010011110";
        when 4824 => y_in <= "10010010"; x_in <= "01011000"; z_correct<="1101101000110000";
        when 4825 => y_in <= "10010010"; x_in <= "01011001"; z_correct<="1101100111000010";
        when 4826 => y_in <= "10010010"; x_in <= "01011010"; z_correct<="1101100101010100";
        when 4827 => y_in <= "10010010"; x_in <= "01011011"; z_correct<="1101100011100110";
        when 4828 => y_in <= "10010010"; x_in <= "01011100"; z_correct<="1101100001111000";
        when 4829 => y_in <= "10010010"; x_in <= "01011101"; z_correct<="1101100000001010";
        when 4830 => y_in <= "10010010"; x_in <= "01011110"; z_correct<="1101011110011100";
        when 4831 => y_in <= "10010010"; x_in <= "01011111"; z_correct<="1101011100101110";
        when 4832 => y_in <= "10010010"; x_in <= "01100000"; z_correct<="1101011011000000";
        when 4833 => y_in <= "10010010"; x_in <= "01100001"; z_correct<="1101011001010010";
        when 4834 => y_in <= "10010010"; x_in <= "01100010"; z_correct<="1101010111100100";
        when 4835 => y_in <= "10010010"; x_in <= "01100011"; z_correct<="1101010101110110";
        when 4836 => y_in <= "10010010"; x_in <= "01100100"; z_correct<="1101010100001000";
        when 4837 => y_in <= "10010010"; x_in <= "01100101"; z_correct<="1101010010011010";
        when 4838 => y_in <= "10010010"; x_in <= "01100110"; z_correct<="1101010000101100";
        when 4839 => y_in <= "10010010"; x_in <= "01100111"; z_correct<="1101001110111110";
        when 4840 => y_in <= "10010010"; x_in <= "01101000"; z_correct<="1101001101010000";
        when 4841 => y_in <= "10010010"; x_in <= "01101001"; z_correct<="1101001011100010";
        when 4842 => y_in <= "10010010"; x_in <= "01101010"; z_correct<="1101001001110100";
        when 4843 => y_in <= "10010010"; x_in <= "01101011"; z_correct<="1101001000000110";
        when 4844 => y_in <= "10010010"; x_in <= "01101100"; z_correct<="1101000110011000";
        when 4845 => y_in <= "10010010"; x_in <= "01101101"; z_correct<="1101000100101010";
        when 4846 => y_in <= "10010010"; x_in <= "01101110"; z_correct<="1101000010111100";
        when 4847 => y_in <= "10010010"; x_in <= "01101111"; z_correct<="1101000001001110";
        when 4848 => y_in <= "10010010"; x_in <= "01110000"; z_correct<="1100111111100000";
        when 4849 => y_in <= "10010010"; x_in <= "01110001"; z_correct<="1100111101110010";
        when 4850 => y_in <= "10010010"; x_in <= "01110010"; z_correct<="1100111100000100";
        when 4851 => y_in <= "10010010"; x_in <= "01110011"; z_correct<="1100111010010110";
        when 4852 => y_in <= "10010010"; x_in <= "01110100"; z_correct<="1100111000101000";
        when 4853 => y_in <= "10010010"; x_in <= "01110101"; z_correct<="1100110110111010";
        when 4854 => y_in <= "10010010"; x_in <= "01110110"; z_correct<="1100110101001100";
        when 4855 => y_in <= "10010010"; x_in <= "01110111"; z_correct<="1100110011011110";
        when 4856 => y_in <= "10010010"; x_in <= "01111000"; z_correct<="1100110001110000";
        when 4857 => y_in <= "10010010"; x_in <= "01111001"; z_correct<="1100110000000010";
        when 4858 => y_in <= "10010010"; x_in <= "01111010"; z_correct<="1100101110010100";
        when 4859 => y_in <= "10010010"; x_in <= "01111011"; z_correct<="1100101100100110";
        when 4860 => y_in <= "10010010"; x_in <= "01111100"; z_correct<="1100101010111000";
        when 4861 => y_in <= "10010010"; x_in <= "01111101"; z_correct<="1100101001001010";
        when 4862 => y_in <= "10010010"; x_in <= "01111110"; z_correct<="1100100111011100";
        when 4863 => y_in <= "10010010"; x_in <= "01111111"; z_correct<="1100100101101110";
        when 4864 => y_in <= "10010011"; x_in <= "10000000"; z_correct<="0011011010000000";
        when 4865 => y_in <= "10010011"; x_in <= "10000001"; z_correct<="0011011000010011";
        when 4866 => y_in <= "10010011"; x_in <= "10000010"; z_correct<="0011010110100110";
        when 4867 => y_in <= "10010011"; x_in <= "10000011"; z_correct<="0011010100111001";
        when 4868 => y_in <= "10010011"; x_in <= "10000100"; z_correct<="0011010011001100";
        when 4869 => y_in <= "10010011"; x_in <= "10000101"; z_correct<="0011010001011111";
        when 4870 => y_in <= "10010011"; x_in <= "10000110"; z_correct<="0011001111110010";
        when 4871 => y_in <= "10010011"; x_in <= "10000111"; z_correct<="0011001110000101";
        when 4872 => y_in <= "10010011"; x_in <= "10001000"; z_correct<="0011001100011000";
        when 4873 => y_in <= "10010011"; x_in <= "10001001"; z_correct<="0011001010101011";
        when 4874 => y_in <= "10010011"; x_in <= "10001010"; z_correct<="0011001000111110";
        when 4875 => y_in <= "10010011"; x_in <= "10001011"; z_correct<="0011000111010001";
        when 4876 => y_in <= "10010011"; x_in <= "10001100"; z_correct<="0011000101100100";
        when 4877 => y_in <= "10010011"; x_in <= "10001101"; z_correct<="0011000011110111";
        when 4878 => y_in <= "10010011"; x_in <= "10001110"; z_correct<="0011000010001010";
        when 4879 => y_in <= "10010011"; x_in <= "10001111"; z_correct<="0011000000011101";
        when 4880 => y_in <= "10010011"; x_in <= "10010000"; z_correct<="0010111110110000";
        when 4881 => y_in <= "10010011"; x_in <= "10010001"; z_correct<="0010111101000011";
        when 4882 => y_in <= "10010011"; x_in <= "10010010"; z_correct<="0010111011010110";
        when 4883 => y_in <= "10010011"; x_in <= "10010011"; z_correct<="0010111001101001";
        when 4884 => y_in <= "10010011"; x_in <= "10010100"; z_correct<="0010110111111100";
        when 4885 => y_in <= "10010011"; x_in <= "10010101"; z_correct<="0010110110001111";
        when 4886 => y_in <= "10010011"; x_in <= "10010110"; z_correct<="0010110100100010";
        when 4887 => y_in <= "10010011"; x_in <= "10010111"; z_correct<="0010110010110101";
        when 4888 => y_in <= "10010011"; x_in <= "10011000"; z_correct<="0010110001001000";
        when 4889 => y_in <= "10010011"; x_in <= "10011001"; z_correct<="0010101111011011";
        when 4890 => y_in <= "10010011"; x_in <= "10011010"; z_correct<="0010101101101110";
        when 4891 => y_in <= "10010011"; x_in <= "10011011"; z_correct<="0010101100000001";
        when 4892 => y_in <= "10010011"; x_in <= "10011100"; z_correct<="0010101010010100";
        when 4893 => y_in <= "10010011"; x_in <= "10011101"; z_correct<="0010101000100111";
        when 4894 => y_in <= "10010011"; x_in <= "10011110"; z_correct<="0010100110111010";
        when 4895 => y_in <= "10010011"; x_in <= "10011111"; z_correct<="0010100101001101";
        when 4896 => y_in <= "10010011"; x_in <= "10100000"; z_correct<="0010100011100000";
        when 4897 => y_in <= "10010011"; x_in <= "10100001"; z_correct<="0010100001110011";
        when 4898 => y_in <= "10010011"; x_in <= "10100010"; z_correct<="0010100000000110";
        when 4899 => y_in <= "10010011"; x_in <= "10100011"; z_correct<="0010011110011001";
        when 4900 => y_in <= "10010011"; x_in <= "10100100"; z_correct<="0010011100101100";
        when 4901 => y_in <= "10010011"; x_in <= "10100101"; z_correct<="0010011010111111";
        when 4902 => y_in <= "10010011"; x_in <= "10100110"; z_correct<="0010011001010010";
        when 4903 => y_in <= "10010011"; x_in <= "10100111"; z_correct<="0010010111100101";
        when 4904 => y_in <= "10010011"; x_in <= "10101000"; z_correct<="0010010101111000";
        when 4905 => y_in <= "10010011"; x_in <= "10101001"; z_correct<="0010010100001011";
        when 4906 => y_in <= "10010011"; x_in <= "10101010"; z_correct<="0010010010011110";
        when 4907 => y_in <= "10010011"; x_in <= "10101011"; z_correct<="0010010000110001";
        when 4908 => y_in <= "10010011"; x_in <= "10101100"; z_correct<="0010001111000100";
        when 4909 => y_in <= "10010011"; x_in <= "10101101"; z_correct<="0010001101010111";
        when 4910 => y_in <= "10010011"; x_in <= "10101110"; z_correct<="0010001011101010";
        when 4911 => y_in <= "10010011"; x_in <= "10101111"; z_correct<="0010001001111101";
        when 4912 => y_in <= "10010011"; x_in <= "10110000"; z_correct<="0010001000010000";
        when 4913 => y_in <= "10010011"; x_in <= "10110001"; z_correct<="0010000110100011";
        when 4914 => y_in <= "10010011"; x_in <= "10110010"; z_correct<="0010000100110110";
        when 4915 => y_in <= "10010011"; x_in <= "10110011"; z_correct<="0010000011001001";
        when 4916 => y_in <= "10010011"; x_in <= "10110100"; z_correct<="0010000001011100";
        when 4917 => y_in <= "10010011"; x_in <= "10110101"; z_correct<="0001111111101111";
        when 4918 => y_in <= "10010011"; x_in <= "10110110"; z_correct<="0001111110000010";
        when 4919 => y_in <= "10010011"; x_in <= "10110111"; z_correct<="0001111100010101";
        when 4920 => y_in <= "10010011"; x_in <= "10111000"; z_correct<="0001111010101000";
        when 4921 => y_in <= "10010011"; x_in <= "10111001"; z_correct<="0001111000111011";
        when 4922 => y_in <= "10010011"; x_in <= "10111010"; z_correct<="0001110111001110";
        when 4923 => y_in <= "10010011"; x_in <= "10111011"; z_correct<="0001110101100001";
        when 4924 => y_in <= "10010011"; x_in <= "10111100"; z_correct<="0001110011110100";
        when 4925 => y_in <= "10010011"; x_in <= "10111101"; z_correct<="0001110010000111";
        when 4926 => y_in <= "10010011"; x_in <= "10111110"; z_correct<="0001110000011010";
        when 4927 => y_in <= "10010011"; x_in <= "10111111"; z_correct<="0001101110101101";
        when 4928 => y_in <= "10010011"; x_in <= "11000000"; z_correct<="0001101101000000";
        when 4929 => y_in <= "10010011"; x_in <= "11000001"; z_correct<="0001101011010011";
        when 4930 => y_in <= "10010011"; x_in <= "11000010"; z_correct<="0001101001100110";
        when 4931 => y_in <= "10010011"; x_in <= "11000011"; z_correct<="0001100111111001";
        when 4932 => y_in <= "10010011"; x_in <= "11000100"; z_correct<="0001100110001100";
        when 4933 => y_in <= "10010011"; x_in <= "11000101"; z_correct<="0001100100011111";
        when 4934 => y_in <= "10010011"; x_in <= "11000110"; z_correct<="0001100010110010";
        when 4935 => y_in <= "10010011"; x_in <= "11000111"; z_correct<="0001100001000101";
        when 4936 => y_in <= "10010011"; x_in <= "11001000"; z_correct<="0001011111011000";
        when 4937 => y_in <= "10010011"; x_in <= "11001001"; z_correct<="0001011101101011";
        when 4938 => y_in <= "10010011"; x_in <= "11001010"; z_correct<="0001011011111110";
        when 4939 => y_in <= "10010011"; x_in <= "11001011"; z_correct<="0001011010010001";
        when 4940 => y_in <= "10010011"; x_in <= "11001100"; z_correct<="0001011000100100";
        when 4941 => y_in <= "10010011"; x_in <= "11001101"; z_correct<="0001010110110111";
        when 4942 => y_in <= "10010011"; x_in <= "11001110"; z_correct<="0001010101001010";
        when 4943 => y_in <= "10010011"; x_in <= "11001111"; z_correct<="0001010011011101";
        when 4944 => y_in <= "10010011"; x_in <= "11010000"; z_correct<="0001010001110000";
        when 4945 => y_in <= "10010011"; x_in <= "11010001"; z_correct<="0001010000000011";
        when 4946 => y_in <= "10010011"; x_in <= "11010010"; z_correct<="0001001110010110";
        when 4947 => y_in <= "10010011"; x_in <= "11010011"; z_correct<="0001001100101001";
        when 4948 => y_in <= "10010011"; x_in <= "11010100"; z_correct<="0001001010111100";
        when 4949 => y_in <= "10010011"; x_in <= "11010101"; z_correct<="0001001001001111";
        when 4950 => y_in <= "10010011"; x_in <= "11010110"; z_correct<="0001000111100010";
        when 4951 => y_in <= "10010011"; x_in <= "11010111"; z_correct<="0001000101110101";
        when 4952 => y_in <= "10010011"; x_in <= "11011000"; z_correct<="0001000100001000";
        when 4953 => y_in <= "10010011"; x_in <= "11011001"; z_correct<="0001000010011011";
        when 4954 => y_in <= "10010011"; x_in <= "11011010"; z_correct<="0001000000101110";
        when 4955 => y_in <= "10010011"; x_in <= "11011011"; z_correct<="0000111111000001";
        when 4956 => y_in <= "10010011"; x_in <= "11011100"; z_correct<="0000111101010100";
        when 4957 => y_in <= "10010011"; x_in <= "11011101"; z_correct<="0000111011100111";
        when 4958 => y_in <= "10010011"; x_in <= "11011110"; z_correct<="0000111001111010";
        when 4959 => y_in <= "10010011"; x_in <= "11011111"; z_correct<="0000111000001101";
        when 4960 => y_in <= "10010011"; x_in <= "11100000"; z_correct<="0000110110100000";
        when 4961 => y_in <= "10010011"; x_in <= "11100001"; z_correct<="0000110100110011";
        when 4962 => y_in <= "10010011"; x_in <= "11100010"; z_correct<="0000110011000110";
        when 4963 => y_in <= "10010011"; x_in <= "11100011"; z_correct<="0000110001011001";
        when 4964 => y_in <= "10010011"; x_in <= "11100100"; z_correct<="0000101111101100";
        when 4965 => y_in <= "10010011"; x_in <= "11100101"; z_correct<="0000101101111111";
        when 4966 => y_in <= "10010011"; x_in <= "11100110"; z_correct<="0000101100010010";
        when 4967 => y_in <= "10010011"; x_in <= "11100111"; z_correct<="0000101010100101";
        when 4968 => y_in <= "10010011"; x_in <= "11101000"; z_correct<="0000101000111000";
        when 4969 => y_in <= "10010011"; x_in <= "11101001"; z_correct<="0000100111001011";
        when 4970 => y_in <= "10010011"; x_in <= "11101010"; z_correct<="0000100101011110";
        when 4971 => y_in <= "10010011"; x_in <= "11101011"; z_correct<="0000100011110001";
        when 4972 => y_in <= "10010011"; x_in <= "11101100"; z_correct<="0000100010000100";
        when 4973 => y_in <= "10010011"; x_in <= "11101101"; z_correct<="0000100000010111";
        when 4974 => y_in <= "10010011"; x_in <= "11101110"; z_correct<="0000011110101010";
        when 4975 => y_in <= "10010011"; x_in <= "11101111"; z_correct<="0000011100111101";
        when 4976 => y_in <= "10010011"; x_in <= "11110000"; z_correct<="0000011011010000";
        when 4977 => y_in <= "10010011"; x_in <= "11110001"; z_correct<="0000011001100011";
        when 4978 => y_in <= "10010011"; x_in <= "11110010"; z_correct<="0000010111110110";
        when 4979 => y_in <= "10010011"; x_in <= "11110011"; z_correct<="0000010110001001";
        when 4980 => y_in <= "10010011"; x_in <= "11110100"; z_correct<="0000010100011100";
        when 4981 => y_in <= "10010011"; x_in <= "11110101"; z_correct<="0000010010101111";
        when 4982 => y_in <= "10010011"; x_in <= "11110110"; z_correct<="0000010001000010";
        when 4983 => y_in <= "10010011"; x_in <= "11110111"; z_correct<="0000001111010101";
        when 4984 => y_in <= "10010011"; x_in <= "11111000"; z_correct<="0000001101101000";
        when 4985 => y_in <= "10010011"; x_in <= "11111001"; z_correct<="0000001011111011";
        when 4986 => y_in <= "10010011"; x_in <= "11111010"; z_correct<="0000001010001110";
        when 4987 => y_in <= "10010011"; x_in <= "11111011"; z_correct<="0000001000100001";
        when 4988 => y_in <= "10010011"; x_in <= "11111100"; z_correct<="0000000110110100";
        when 4989 => y_in <= "10010011"; x_in <= "11111101"; z_correct<="0000000101000111";
        when 4990 => y_in <= "10010011"; x_in <= "11111110"; z_correct<="0000000011011010";
        when 4991 => y_in <= "10010011"; x_in <= "11111111"; z_correct<="0000000001101101";
        when 4992 => y_in <= "10010011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 4993 => y_in <= "10010011"; x_in <= "00000001"; z_correct<="1111111110010011";
        when 4994 => y_in <= "10010011"; x_in <= "00000010"; z_correct<="1111111100100110";
        when 4995 => y_in <= "10010011"; x_in <= "00000011"; z_correct<="1111111010111001";
        when 4996 => y_in <= "10010011"; x_in <= "00000100"; z_correct<="1111111001001100";
        when 4997 => y_in <= "10010011"; x_in <= "00000101"; z_correct<="1111110111011111";
        when 4998 => y_in <= "10010011"; x_in <= "00000110"; z_correct<="1111110101110010";
        when 4999 => y_in <= "10010011"; x_in <= "00000111"; z_correct<="1111110100000101";
        when 5000 => y_in <= "10010011"; x_in <= "00001000"; z_correct<="1111110010011000";
        when 5001 => y_in <= "10010011"; x_in <= "00001001"; z_correct<="1111110000101011";
        when 5002 => y_in <= "10010011"; x_in <= "00001010"; z_correct<="1111101110111110";
        when 5003 => y_in <= "10010011"; x_in <= "00001011"; z_correct<="1111101101010001";
        when 5004 => y_in <= "10010011"; x_in <= "00001100"; z_correct<="1111101011100100";
        when 5005 => y_in <= "10010011"; x_in <= "00001101"; z_correct<="1111101001110111";
        when 5006 => y_in <= "10010011"; x_in <= "00001110"; z_correct<="1111101000001010";
        when 5007 => y_in <= "10010011"; x_in <= "00001111"; z_correct<="1111100110011101";
        when 5008 => y_in <= "10010011"; x_in <= "00010000"; z_correct<="1111100100110000";
        when 5009 => y_in <= "10010011"; x_in <= "00010001"; z_correct<="1111100011000011";
        when 5010 => y_in <= "10010011"; x_in <= "00010010"; z_correct<="1111100001010110";
        when 5011 => y_in <= "10010011"; x_in <= "00010011"; z_correct<="1111011111101001";
        when 5012 => y_in <= "10010011"; x_in <= "00010100"; z_correct<="1111011101111100";
        when 5013 => y_in <= "10010011"; x_in <= "00010101"; z_correct<="1111011100001111";
        when 5014 => y_in <= "10010011"; x_in <= "00010110"; z_correct<="1111011010100010";
        when 5015 => y_in <= "10010011"; x_in <= "00010111"; z_correct<="1111011000110101";
        when 5016 => y_in <= "10010011"; x_in <= "00011000"; z_correct<="1111010111001000";
        when 5017 => y_in <= "10010011"; x_in <= "00011001"; z_correct<="1111010101011011";
        when 5018 => y_in <= "10010011"; x_in <= "00011010"; z_correct<="1111010011101110";
        when 5019 => y_in <= "10010011"; x_in <= "00011011"; z_correct<="1111010010000001";
        when 5020 => y_in <= "10010011"; x_in <= "00011100"; z_correct<="1111010000010100";
        when 5021 => y_in <= "10010011"; x_in <= "00011101"; z_correct<="1111001110100111";
        when 5022 => y_in <= "10010011"; x_in <= "00011110"; z_correct<="1111001100111010";
        when 5023 => y_in <= "10010011"; x_in <= "00011111"; z_correct<="1111001011001101";
        when 5024 => y_in <= "10010011"; x_in <= "00100000"; z_correct<="1111001001100000";
        when 5025 => y_in <= "10010011"; x_in <= "00100001"; z_correct<="1111000111110011";
        when 5026 => y_in <= "10010011"; x_in <= "00100010"; z_correct<="1111000110000110";
        when 5027 => y_in <= "10010011"; x_in <= "00100011"; z_correct<="1111000100011001";
        when 5028 => y_in <= "10010011"; x_in <= "00100100"; z_correct<="1111000010101100";
        when 5029 => y_in <= "10010011"; x_in <= "00100101"; z_correct<="1111000000111111";
        when 5030 => y_in <= "10010011"; x_in <= "00100110"; z_correct<="1110111111010010";
        when 5031 => y_in <= "10010011"; x_in <= "00100111"; z_correct<="1110111101100101";
        when 5032 => y_in <= "10010011"; x_in <= "00101000"; z_correct<="1110111011111000";
        when 5033 => y_in <= "10010011"; x_in <= "00101001"; z_correct<="1110111010001011";
        when 5034 => y_in <= "10010011"; x_in <= "00101010"; z_correct<="1110111000011110";
        when 5035 => y_in <= "10010011"; x_in <= "00101011"; z_correct<="1110110110110001";
        when 5036 => y_in <= "10010011"; x_in <= "00101100"; z_correct<="1110110101000100";
        when 5037 => y_in <= "10010011"; x_in <= "00101101"; z_correct<="1110110011010111";
        when 5038 => y_in <= "10010011"; x_in <= "00101110"; z_correct<="1110110001101010";
        when 5039 => y_in <= "10010011"; x_in <= "00101111"; z_correct<="1110101111111101";
        when 5040 => y_in <= "10010011"; x_in <= "00110000"; z_correct<="1110101110010000";
        when 5041 => y_in <= "10010011"; x_in <= "00110001"; z_correct<="1110101100100011";
        when 5042 => y_in <= "10010011"; x_in <= "00110010"; z_correct<="1110101010110110";
        when 5043 => y_in <= "10010011"; x_in <= "00110011"; z_correct<="1110101001001001";
        when 5044 => y_in <= "10010011"; x_in <= "00110100"; z_correct<="1110100111011100";
        when 5045 => y_in <= "10010011"; x_in <= "00110101"; z_correct<="1110100101101111";
        when 5046 => y_in <= "10010011"; x_in <= "00110110"; z_correct<="1110100100000010";
        when 5047 => y_in <= "10010011"; x_in <= "00110111"; z_correct<="1110100010010101";
        when 5048 => y_in <= "10010011"; x_in <= "00111000"; z_correct<="1110100000101000";
        when 5049 => y_in <= "10010011"; x_in <= "00111001"; z_correct<="1110011110111011";
        when 5050 => y_in <= "10010011"; x_in <= "00111010"; z_correct<="1110011101001110";
        when 5051 => y_in <= "10010011"; x_in <= "00111011"; z_correct<="1110011011100001";
        when 5052 => y_in <= "10010011"; x_in <= "00111100"; z_correct<="1110011001110100";
        when 5053 => y_in <= "10010011"; x_in <= "00111101"; z_correct<="1110011000000111";
        when 5054 => y_in <= "10010011"; x_in <= "00111110"; z_correct<="1110010110011010";
        when 5055 => y_in <= "10010011"; x_in <= "00111111"; z_correct<="1110010100101101";
        when 5056 => y_in <= "10010011"; x_in <= "01000000"; z_correct<="1110010011000000";
        when 5057 => y_in <= "10010011"; x_in <= "01000001"; z_correct<="1110010001010011";
        when 5058 => y_in <= "10010011"; x_in <= "01000010"; z_correct<="1110001111100110";
        when 5059 => y_in <= "10010011"; x_in <= "01000011"; z_correct<="1110001101111001";
        when 5060 => y_in <= "10010011"; x_in <= "01000100"; z_correct<="1110001100001100";
        when 5061 => y_in <= "10010011"; x_in <= "01000101"; z_correct<="1110001010011111";
        when 5062 => y_in <= "10010011"; x_in <= "01000110"; z_correct<="1110001000110010";
        when 5063 => y_in <= "10010011"; x_in <= "01000111"; z_correct<="1110000111000101";
        when 5064 => y_in <= "10010011"; x_in <= "01001000"; z_correct<="1110000101011000";
        when 5065 => y_in <= "10010011"; x_in <= "01001001"; z_correct<="1110000011101011";
        when 5066 => y_in <= "10010011"; x_in <= "01001010"; z_correct<="1110000001111110";
        when 5067 => y_in <= "10010011"; x_in <= "01001011"; z_correct<="1110000000010001";
        when 5068 => y_in <= "10010011"; x_in <= "01001100"; z_correct<="1101111110100100";
        when 5069 => y_in <= "10010011"; x_in <= "01001101"; z_correct<="1101111100110111";
        when 5070 => y_in <= "10010011"; x_in <= "01001110"; z_correct<="1101111011001010";
        when 5071 => y_in <= "10010011"; x_in <= "01001111"; z_correct<="1101111001011101";
        when 5072 => y_in <= "10010011"; x_in <= "01010000"; z_correct<="1101110111110000";
        when 5073 => y_in <= "10010011"; x_in <= "01010001"; z_correct<="1101110110000011";
        when 5074 => y_in <= "10010011"; x_in <= "01010010"; z_correct<="1101110100010110";
        when 5075 => y_in <= "10010011"; x_in <= "01010011"; z_correct<="1101110010101001";
        when 5076 => y_in <= "10010011"; x_in <= "01010100"; z_correct<="1101110000111100";
        when 5077 => y_in <= "10010011"; x_in <= "01010101"; z_correct<="1101101111001111";
        when 5078 => y_in <= "10010011"; x_in <= "01010110"; z_correct<="1101101101100010";
        when 5079 => y_in <= "10010011"; x_in <= "01010111"; z_correct<="1101101011110101";
        when 5080 => y_in <= "10010011"; x_in <= "01011000"; z_correct<="1101101010001000";
        when 5081 => y_in <= "10010011"; x_in <= "01011001"; z_correct<="1101101000011011";
        when 5082 => y_in <= "10010011"; x_in <= "01011010"; z_correct<="1101100110101110";
        when 5083 => y_in <= "10010011"; x_in <= "01011011"; z_correct<="1101100101000001";
        when 5084 => y_in <= "10010011"; x_in <= "01011100"; z_correct<="1101100011010100";
        when 5085 => y_in <= "10010011"; x_in <= "01011101"; z_correct<="1101100001100111";
        when 5086 => y_in <= "10010011"; x_in <= "01011110"; z_correct<="1101011111111010";
        when 5087 => y_in <= "10010011"; x_in <= "01011111"; z_correct<="1101011110001101";
        when 5088 => y_in <= "10010011"; x_in <= "01100000"; z_correct<="1101011100100000";
        when 5089 => y_in <= "10010011"; x_in <= "01100001"; z_correct<="1101011010110011";
        when 5090 => y_in <= "10010011"; x_in <= "01100010"; z_correct<="1101011001000110";
        when 5091 => y_in <= "10010011"; x_in <= "01100011"; z_correct<="1101010111011001";
        when 5092 => y_in <= "10010011"; x_in <= "01100100"; z_correct<="1101010101101100";
        when 5093 => y_in <= "10010011"; x_in <= "01100101"; z_correct<="1101010011111111";
        when 5094 => y_in <= "10010011"; x_in <= "01100110"; z_correct<="1101010010010010";
        when 5095 => y_in <= "10010011"; x_in <= "01100111"; z_correct<="1101010000100101";
        when 5096 => y_in <= "10010011"; x_in <= "01101000"; z_correct<="1101001110111000";
        when 5097 => y_in <= "10010011"; x_in <= "01101001"; z_correct<="1101001101001011";
        when 5098 => y_in <= "10010011"; x_in <= "01101010"; z_correct<="1101001011011110";
        when 5099 => y_in <= "10010011"; x_in <= "01101011"; z_correct<="1101001001110001";
        when 5100 => y_in <= "10010011"; x_in <= "01101100"; z_correct<="1101001000000100";
        when 5101 => y_in <= "10010011"; x_in <= "01101101"; z_correct<="1101000110010111";
        when 5102 => y_in <= "10010011"; x_in <= "01101110"; z_correct<="1101000100101010";
        when 5103 => y_in <= "10010011"; x_in <= "01101111"; z_correct<="1101000010111101";
        when 5104 => y_in <= "10010011"; x_in <= "01110000"; z_correct<="1101000001010000";
        when 5105 => y_in <= "10010011"; x_in <= "01110001"; z_correct<="1100111111100011";
        when 5106 => y_in <= "10010011"; x_in <= "01110010"; z_correct<="1100111101110110";
        when 5107 => y_in <= "10010011"; x_in <= "01110011"; z_correct<="1100111100001001";
        when 5108 => y_in <= "10010011"; x_in <= "01110100"; z_correct<="1100111010011100";
        when 5109 => y_in <= "10010011"; x_in <= "01110101"; z_correct<="1100111000101111";
        when 5110 => y_in <= "10010011"; x_in <= "01110110"; z_correct<="1100110111000010";
        when 5111 => y_in <= "10010011"; x_in <= "01110111"; z_correct<="1100110101010101";
        when 5112 => y_in <= "10010011"; x_in <= "01111000"; z_correct<="1100110011101000";
        when 5113 => y_in <= "10010011"; x_in <= "01111001"; z_correct<="1100110001111011";
        when 5114 => y_in <= "10010011"; x_in <= "01111010"; z_correct<="1100110000001110";
        when 5115 => y_in <= "10010011"; x_in <= "01111011"; z_correct<="1100101110100001";
        when 5116 => y_in <= "10010011"; x_in <= "01111100"; z_correct<="1100101100110100";
        when 5117 => y_in <= "10010011"; x_in <= "01111101"; z_correct<="1100101011000111";
        when 5118 => y_in <= "10010011"; x_in <= "01111110"; z_correct<="1100101001011010";
        when 5119 => y_in <= "10010011"; x_in <= "01111111"; z_correct<="1100100111101101";
        when 5120 => y_in <= "10010100"; x_in <= "10000000"; z_correct<="0011011000000000";
        when 5121 => y_in <= "10010100"; x_in <= "10000001"; z_correct<="0011010110010100";
        when 5122 => y_in <= "10010100"; x_in <= "10000010"; z_correct<="0011010100101000";
        when 5123 => y_in <= "10010100"; x_in <= "10000011"; z_correct<="0011010010111100";
        when 5124 => y_in <= "10010100"; x_in <= "10000100"; z_correct<="0011010001010000";
        when 5125 => y_in <= "10010100"; x_in <= "10000101"; z_correct<="0011001111100100";
        when 5126 => y_in <= "10010100"; x_in <= "10000110"; z_correct<="0011001101111000";
        when 5127 => y_in <= "10010100"; x_in <= "10000111"; z_correct<="0011001100001100";
        when 5128 => y_in <= "10010100"; x_in <= "10001000"; z_correct<="0011001010100000";
        when 5129 => y_in <= "10010100"; x_in <= "10001001"; z_correct<="0011001000110100";
        when 5130 => y_in <= "10010100"; x_in <= "10001010"; z_correct<="0011000111001000";
        when 5131 => y_in <= "10010100"; x_in <= "10001011"; z_correct<="0011000101011100";
        when 5132 => y_in <= "10010100"; x_in <= "10001100"; z_correct<="0011000011110000";
        when 5133 => y_in <= "10010100"; x_in <= "10001101"; z_correct<="0011000010000100";
        when 5134 => y_in <= "10010100"; x_in <= "10001110"; z_correct<="0011000000011000";
        when 5135 => y_in <= "10010100"; x_in <= "10001111"; z_correct<="0010111110101100";
        when 5136 => y_in <= "10010100"; x_in <= "10010000"; z_correct<="0010111101000000";
        when 5137 => y_in <= "10010100"; x_in <= "10010001"; z_correct<="0010111011010100";
        when 5138 => y_in <= "10010100"; x_in <= "10010010"; z_correct<="0010111001101000";
        when 5139 => y_in <= "10010100"; x_in <= "10010011"; z_correct<="0010110111111100";
        when 5140 => y_in <= "10010100"; x_in <= "10010100"; z_correct<="0010110110010000";
        when 5141 => y_in <= "10010100"; x_in <= "10010101"; z_correct<="0010110100100100";
        when 5142 => y_in <= "10010100"; x_in <= "10010110"; z_correct<="0010110010111000";
        when 5143 => y_in <= "10010100"; x_in <= "10010111"; z_correct<="0010110001001100";
        when 5144 => y_in <= "10010100"; x_in <= "10011000"; z_correct<="0010101111100000";
        when 5145 => y_in <= "10010100"; x_in <= "10011001"; z_correct<="0010101101110100";
        when 5146 => y_in <= "10010100"; x_in <= "10011010"; z_correct<="0010101100001000";
        when 5147 => y_in <= "10010100"; x_in <= "10011011"; z_correct<="0010101010011100";
        when 5148 => y_in <= "10010100"; x_in <= "10011100"; z_correct<="0010101000110000";
        when 5149 => y_in <= "10010100"; x_in <= "10011101"; z_correct<="0010100111000100";
        when 5150 => y_in <= "10010100"; x_in <= "10011110"; z_correct<="0010100101011000";
        when 5151 => y_in <= "10010100"; x_in <= "10011111"; z_correct<="0010100011101100";
        when 5152 => y_in <= "10010100"; x_in <= "10100000"; z_correct<="0010100010000000";
        when 5153 => y_in <= "10010100"; x_in <= "10100001"; z_correct<="0010100000010100";
        when 5154 => y_in <= "10010100"; x_in <= "10100010"; z_correct<="0010011110101000";
        when 5155 => y_in <= "10010100"; x_in <= "10100011"; z_correct<="0010011100111100";
        when 5156 => y_in <= "10010100"; x_in <= "10100100"; z_correct<="0010011011010000";
        when 5157 => y_in <= "10010100"; x_in <= "10100101"; z_correct<="0010011001100100";
        when 5158 => y_in <= "10010100"; x_in <= "10100110"; z_correct<="0010010111111000";
        when 5159 => y_in <= "10010100"; x_in <= "10100111"; z_correct<="0010010110001100";
        when 5160 => y_in <= "10010100"; x_in <= "10101000"; z_correct<="0010010100100000";
        when 5161 => y_in <= "10010100"; x_in <= "10101001"; z_correct<="0010010010110100";
        when 5162 => y_in <= "10010100"; x_in <= "10101010"; z_correct<="0010010001001000";
        when 5163 => y_in <= "10010100"; x_in <= "10101011"; z_correct<="0010001111011100";
        when 5164 => y_in <= "10010100"; x_in <= "10101100"; z_correct<="0010001101110000";
        when 5165 => y_in <= "10010100"; x_in <= "10101101"; z_correct<="0010001100000100";
        when 5166 => y_in <= "10010100"; x_in <= "10101110"; z_correct<="0010001010011000";
        when 5167 => y_in <= "10010100"; x_in <= "10101111"; z_correct<="0010001000101100";
        when 5168 => y_in <= "10010100"; x_in <= "10110000"; z_correct<="0010000111000000";
        when 5169 => y_in <= "10010100"; x_in <= "10110001"; z_correct<="0010000101010100";
        when 5170 => y_in <= "10010100"; x_in <= "10110010"; z_correct<="0010000011101000";
        when 5171 => y_in <= "10010100"; x_in <= "10110011"; z_correct<="0010000001111100";
        when 5172 => y_in <= "10010100"; x_in <= "10110100"; z_correct<="0010000000010000";
        when 5173 => y_in <= "10010100"; x_in <= "10110101"; z_correct<="0001111110100100";
        when 5174 => y_in <= "10010100"; x_in <= "10110110"; z_correct<="0001111100111000";
        when 5175 => y_in <= "10010100"; x_in <= "10110111"; z_correct<="0001111011001100";
        when 5176 => y_in <= "10010100"; x_in <= "10111000"; z_correct<="0001111001100000";
        when 5177 => y_in <= "10010100"; x_in <= "10111001"; z_correct<="0001110111110100";
        when 5178 => y_in <= "10010100"; x_in <= "10111010"; z_correct<="0001110110001000";
        when 5179 => y_in <= "10010100"; x_in <= "10111011"; z_correct<="0001110100011100";
        when 5180 => y_in <= "10010100"; x_in <= "10111100"; z_correct<="0001110010110000";
        when 5181 => y_in <= "10010100"; x_in <= "10111101"; z_correct<="0001110001000100";
        when 5182 => y_in <= "10010100"; x_in <= "10111110"; z_correct<="0001101111011000";
        when 5183 => y_in <= "10010100"; x_in <= "10111111"; z_correct<="0001101101101100";
        when 5184 => y_in <= "10010100"; x_in <= "11000000"; z_correct<="0001101100000000";
        when 5185 => y_in <= "10010100"; x_in <= "11000001"; z_correct<="0001101010010100";
        when 5186 => y_in <= "10010100"; x_in <= "11000010"; z_correct<="0001101000101000";
        when 5187 => y_in <= "10010100"; x_in <= "11000011"; z_correct<="0001100110111100";
        when 5188 => y_in <= "10010100"; x_in <= "11000100"; z_correct<="0001100101010000";
        when 5189 => y_in <= "10010100"; x_in <= "11000101"; z_correct<="0001100011100100";
        when 5190 => y_in <= "10010100"; x_in <= "11000110"; z_correct<="0001100001111000";
        when 5191 => y_in <= "10010100"; x_in <= "11000111"; z_correct<="0001100000001100";
        when 5192 => y_in <= "10010100"; x_in <= "11001000"; z_correct<="0001011110100000";
        when 5193 => y_in <= "10010100"; x_in <= "11001001"; z_correct<="0001011100110100";
        when 5194 => y_in <= "10010100"; x_in <= "11001010"; z_correct<="0001011011001000";
        when 5195 => y_in <= "10010100"; x_in <= "11001011"; z_correct<="0001011001011100";
        when 5196 => y_in <= "10010100"; x_in <= "11001100"; z_correct<="0001010111110000";
        when 5197 => y_in <= "10010100"; x_in <= "11001101"; z_correct<="0001010110000100";
        when 5198 => y_in <= "10010100"; x_in <= "11001110"; z_correct<="0001010100011000";
        when 5199 => y_in <= "10010100"; x_in <= "11001111"; z_correct<="0001010010101100";
        when 5200 => y_in <= "10010100"; x_in <= "11010000"; z_correct<="0001010001000000";
        when 5201 => y_in <= "10010100"; x_in <= "11010001"; z_correct<="0001001111010100";
        when 5202 => y_in <= "10010100"; x_in <= "11010010"; z_correct<="0001001101101000";
        when 5203 => y_in <= "10010100"; x_in <= "11010011"; z_correct<="0001001011111100";
        when 5204 => y_in <= "10010100"; x_in <= "11010100"; z_correct<="0001001010010000";
        when 5205 => y_in <= "10010100"; x_in <= "11010101"; z_correct<="0001001000100100";
        when 5206 => y_in <= "10010100"; x_in <= "11010110"; z_correct<="0001000110111000";
        when 5207 => y_in <= "10010100"; x_in <= "11010111"; z_correct<="0001000101001100";
        when 5208 => y_in <= "10010100"; x_in <= "11011000"; z_correct<="0001000011100000";
        when 5209 => y_in <= "10010100"; x_in <= "11011001"; z_correct<="0001000001110100";
        when 5210 => y_in <= "10010100"; x_in <= "11011010"; z_correct<="0001000000001000";
        when 5211 => y_in <= "10010100"; x_in <= "11011011"; z_correct<="0000111110011100";
        when 5212 => y_in <= "10010100"; x_in <= "11011100"; z_correct<="0000111100110000";
        when 5213 => y_in <= "10010100"; x_in <= "11011101"; z_correct<="0000111011000100";
        when 5214 => y_in <= "10010100"; x_in <= "11011110"; z_correct<="0000111001011000";
        when 5215 => y_in <= "10010100"; x_in <= "11011111"; z_correct<="0000110111101100";
        when 5216 => y_in <= "10010100"; x_in <= "11100000"; z_correct<="0000110110000000";
        when 5217 => y_in <= "10010100"; x_in <= "11100001"; z_correct<="0000110100010100";
        when 5218 => y_in <= "10010100"; x_in <= "11100010"; z_correct<="0000110010101000";
        when 5219 => y_in <= "10010100"; x_in <= "11100011"; z_correct<="0000110000111100";
        when 5220 => y_in <= "10010100"; x_in <= "11100100"; z_correct<="0000101111010000";
        when 5221 => y_in <= "10010100"; x_in <= "11100101"; z_correct<="0000101101100100";
        when 5222 => y_in <= "10010100"; x_in <= "11100110"; z_correct<="0000101011111000";
        when 5223 => y_in <= "10010100"; x_in <= "11100111"; z_correct<="0000101010001100";
        when 5224 => y_in <= "10010100"; x_in <= "11101000"; z_correct<="0000101000100000";
        when 5225 => y_in <= "10010100"; x_in <= "11101001"; z_correct<="0000100110110100";
        when 5226 => y_in <= "10010100"; x_in <= "11101010"; z_correct<="0000100101001000";
        when 5227 => y_in <= "10010100"; x_in <= "11101011"; z_correct<="0000100011011100";
        when 5228 => y_in <= "10010100"; x_in <= "11101100"; z_correct<="0000100001110000";
        when 5229 => y_in <= "10010100"; x_in <= "11101101"; z_correct<="0000100000000100";
        when 5230 => y_in <= "10010100"; x_in <= "11101110"; z_correct<="0000011110011000";
        when 5231 => y_in <= "10010100"; x_in <= "11101111"; z_correct<="0000011100101100";
        when 5232 => y_in <= "10010100"; x_in <= "11110000"; z_correct<="0000011011000000";
        when 5233 => y_in <= "10010100"; x_in <= "11110001"; z_correct<="0000011001010100";
        when 5234 => y_in <= "10010100"; x_in <= "11110010"; z_correct<="0000010111101000";
        when 5235 => y_in <= "10010100"; x_in <= "11110011"; z_correct<="0000010101111100";
        when 5236 => y_in <= "10010100"; x_in <= "11110100"; z_correct<="0000010100010000";
        when 5237 => y_in <= "10010100"; x_in <= "11110101"; z_correct<="0000010010100100";
        when 5238 => y_in <= "10010100"; x_in <= "11110110"; z_correct<="0000010000111000";
        when 5239 => y_in <= "10010100"; x_in <= "11110111"; z_correct<="0000001111001100";
        when 5240 => y_in <= "10010100"; x_in <= "11111000"; z_correct<="0000001101100000";
        when 5241 => y_in <= "10010100"; x_in <= "11111001"; z_correct<="0000001011110100";
        when 5242 => y_in <= "10010100"; x_in <= "11111010"; z_correct<="0000001010001000";
        when 5243 => y_in <= "10010100"; x_in <= "11111011"; z_correct<="0000001000011100";
        when 5244 => y_in <= "10010100"; x_in <= "11111100"; z_correct<="0000000110110000";
        when 5245 => y_in <= "10010100"; x_in <= "11111101"; z_correct<="0000000101000100";
        when 5246 => y_in <= "10010100"; x_in <= "11111110"; z_correct<="0000000011011000";
        when 5247 => y_in <= "10010100"; x_in <= "11111111"; z_correct<="0000000001101100";
        when 5248 => y_in <= "10010100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 5249 => y_in <= "10010100"; x_in <= "00000001"; z_correct<="1111111110010100";
        when 5250 => y_in <= "10010100"; x_in <= "00000010"; z_correct<="1111111100101000";
        when 5251 => y_in <= "10010100"; x_in <= "00000011"; z_correct<="1111111010111100";
        when 5252 => y_in <= "10010100"; x_in <= "00000100"; z_correct<="1111111001010000";
        when 5253 => y_in <= "10010100"; x_in <= "00000101"; z_correct<="1111110111100100";
        when 5254 => y_in <= "10010100"; x_in <= "00000110"; z_correct<="1111110101111000";
        when 5255 => y_in <= "10010100"; x_in <= "00000111"; z_correct<="1111110100001100";
        when 5256 => y_in <= "10010100"; x_in <= "00001000"; z_correct<="1111110010100000";
        when 5257 => y_in <= "10010100"; x_in <= "00001001"; z_correct<="1111110000110100";
        when 5258 => y_in <= "10010100"; x_in <= "00001010"; z_correct<="1111101111001000";
        when 5259 => y_in <= "10010100"; x_in <= "00001011"; z_correct<="1111101101011100";
        when 5260 => y_in <= "10010100"; x_in <= "00001100"; z_correct<="1111101011110000";
        when 5261 => y_in <= "10010100"; x_in <= "00001101"; z_correct<="1111101010000100";
        when 5262 => y_in <= "10010100"; x_in <= "00001110"; z_correct<="1111101000011000";
        when 5263 => y_in <= "10010100"; x_in <= "00001111"; z_correct<="1111100110101100";
        when 5264 => y_in <= "10010100"; x_in <= "00010000"; z_correct<="1111100101000000";
        when 5265 => y_in <= "10010100"; x_in <= "00010001"; z_correct<="1111100011010100";
        when 5266 => y_in <= "10010100"; x_in <= "00010010"; z_correct<="1111100001101000";
        when 5267 => y_in <= "10010100"; x_in <= "00010011"; z_correct<="1111011111111100";
        when 5268 => y_in <= "10010100"; x_in <= "00010100"; z_correct<="1111011110010000";
        when 5269 => y_in <= "10010100"; x_in <= "00010101"; z_correct<="1111011100100100";
        when 5270 => y_in <= "10010100"; x_in <= "00010110"; z_correct<="1111011010111000";
        when 5271 => y_in <= "10010100"; x_in <= "00010111"; z_correct<="1111011001001100";
        when 5272 => y_in <= "10010100"; x_in <= "00011000"; z_correct<="1111010111100000";
        when 5273 => y_in <= "10010100"; x_in <= "00011001"; z_correct<="1111010101110100";
        when 5274 => y_in <= "10010100"; x_in <= "00011010"; z_correct<="1111010100001000";
        when 5275 => y_in <= "10010100"; x_in <= "00011011"; z_correct<="1111010010011100";
        when 5276 => y_in <= "10010100"; x_in <= "00011100"; z_correct<="1111010000110000";
        when 5277 => y_in <= "10010100"; x_in <= "00011101"; z_correct<="1111001111000100";
        when 5278 => y_in <= "10010100"; x_in <= "00011110"; z_correct<="1111001101011000";
        when 5279 => y_in <= "10010100"; x_in <= "00011111"; z_correct<="1111001011101100";
        when 5280 => y_in <= "10010100"; x_in <= "00100000"; z_correct<="1111001010000000";
        when 5281 => y_in <= "10010100"; x_in <= "00100001"; z_correct<="1111001000010100";
        when 5282 => y_in <= "10010100"; x_in <= "00100010"; z_correct<="1111000110101000";
        when 5283 => y_in <= "10010100"; x_in <= "00100011"; z_correct<="1111000100111100";
        when 5284 => y_in <= "10010100"; x_in <= "00100100"; z_correct<="1111000011010000";
        when 5285 => y_in <= "10010100"; x_in <= "00100101"; z_correct<="1111000001100100";
        when 5286 => y_in <= "10010100"; x_in <= "00100110"; z_correct<="1110111111111000";
        when 5287 => y_in <= "10010100"; x_in <= "00100111"; z_correct<="1110111110001100";
        when 5288 => y_in <= "10010100"; x_in <= "00101000"; z_correct<="1110111100100000";
        when 5289 => y_in <= "10010100"; x_in <= "00101001"; z_correct<="1110111010110100";
        when 5290 => y_in <= "10010100"; x_in <= "00101010"; z_correct<="1110111001001000";
        when 5291 => y_in <= "10010100"; x_in <= "00101011"; z_correct<="1110110111011100";
        when 5292 => y_in <= "10010100"; x_in <= "00101100"; z_correct<="1110110101110000";
        when 5293 => y_in <= "10010100"; x_in <= "00101101"; z_correct<="1110110100000100";
        when 5294 => y_in <= "10010100"; x_in <= "00101110"; z_correct<="1110110010011000";
        when 5295 => y_in <= "10010100"; x_in <= "00101111"; z_correct<="1110110000101100";
        when 5296 => y_in <= "10010100"; x_in <= "00110000"; z_correct<="1110101111000000";
        when 5297 => y_in <= "10010100"; x_in <= "00110001"; z_correct<="1110101101010100";
        when 5298 => y_in <= "10010100"; x_in <= "00110010"; z_correct<="1110101011101000";
        when 5299 => y_in <= "10010100"; x_in <= "00110011"; z_correct<="1110101001111100";
        when 5300 => y_in <= "10010100"; x_in <= "00110100"; z_correct<="1110101000010000";
        when 5301 => y_in <= "10010100"; x_in <= "00110101"; z_correct<="1110100110100100";
        when 5302 => y_in <= "10010100"; x_in <= "00110110"; z_correct<="1110100100111000";
        when 5303 => y_in <= "10010100"; x_in <= "00110111"; z_correct<="1110100011001100";
        when 5304 => y_in <= "10010100"; x_in <= "00111000"; z_correct<="1110100001100000";
        when 5305 => y_in <= "10010100"; x_in <= "00111001"; z_correct<="1110011111110100";
        when 5306 => y_in <= "10010100"; x_in <= "00111010"; z_correct<="1110011110001000";
        when 5307 => y_in <= "10010100"; x_in <= "00111011"; z_correct<="1110011100011100";
        when 5308 => y_in <= "10010100"; x_in <= "00111100"; z_correct<="1110011010110000";
        when 5309 => y_in <= "10010100"; x_in <= "00111101"; z_correct<="1110011001000100";
        when 5310 => y_in <= "10010100"; x_in <= "00111110"; z_correct<="1110010111011000";
        when 5311 => y_in <= "10010100"; x_in <= "00111111"; z_correct<="1110010101101100";
        when 5312 => y_in <= "10010100"; x_in <= "01000000"; z_correct<="1110010100000000";
        when 5313 => y_in <= "10010100"; x_in <= "01000001"; z_correct<="1110010010010100";
        when 5314 => y_in <= "10010100"; x_in <= "01000010"; z_correct<="1110010000101000";
        when 5315 => y_in <= "10010100"; x_in <= "01000011"; z_correct<="1110001110111100";
        when 5316 => y_in <= "10010100"; x_in <= "01000100"; z_correct<="1110001101010000";
        when 5317 => y_in <= "10010100"; x_in <= "01000101"; z_correct<="1110001011100100";
        when 5318 => y_in <= "10010100"; x_in <= "01000110"; z_correct<="1110001001111000";
        when 5319 => y_in <= "10010100"; x_in <= "01000111"; z_correct<="1110001000001100";
        when 5320 => y_in <= "10010100"; x_in <= "01001000"; z_correct<="1110000110100000";
        when 5321 => y_in <= "10010100"; x_in <= "01001001"; z_correct<="1110000100110100";
        when 5322 => y_in <= "10010100"; x_in <= "01001010"; z_correct<="1110000011001000";
        when 5323 => y_in <= "10010100"; x_in <= "01001011"; z_correct<="1110000001011100";
        when 5324 => y_in <= "10010100"; x_in <= "01001100"; z_correct<="1101111111110000";
        when 5325 => y_in <= "10010100"; x_in <= "01001101"; z_correct<="1101111110000100";
        when 5326 => y_in <= "10010100"; x_in <= "01001110"; z_correct<="1101111100011000";
        when 5327 => y_in <= "10010100"; x_in <= "01001111"; z_correct<="1101111010101100";
        when 5328 => y_in <= "10010100"; x_in <= "01010000"; z_correct<="1101111001000000";
        when 5329 => y_in <= "10010100"; x_in <= "01010001"; z_correct<="1101110111010100";
        when 5330 => y_in <= "10010100"; x_in <= "01010010"; z_correct<="1101110101101000";
        when 5331 => y_in <= "10010100"; x_in <= "01010011"; z_correct<="1101110011111100";
        when 5332 => y_in <= "10010100"; x_in <= "01010100"; z_correct<="1101110010010000";
        when 5333 => y_in <= "10010100"; x_in <= "01010101"; z_correct<="1101110000100100";
        when 5334 => y_in <= "10010100"; x_in <= "01010110"; z_correct<="1101101110111000";
        when 5335 => y_in <= "10010100"; x_in <= "01010111"; z_correct<="1101101101001100";
        when 5336 => y_in <= "10010100"; x_in <= "01011000"; z_correct<="1101101011100000";
        when 5337 => y_in <= "10010100"; x_in <= "01011001"; z_correct<="1101101001110100";
        when 5338 => y_in <= "10010100"; x_in <= "01011010"; z_correct<="1101101000001000";
        when 5339 => y_in <= "10010100"; x_in <= "01011011"; z_correct<="1101100110011100";
        when 5340 => y_in <= "10010100"; x_in <= "01011100"; z_correct<="1101100100110000";
        when 5341 => y_in <= "10010100"; x_in <= "01011101"; z_correct<="1101100011000100";
        when 5342 => y_in <= "10010100"; x_in <= "01011110"; z_correct<="1101100001011000";
        when 5343 => y_in <= "10010100"; x_in <= "01011111"; z_correct<="1101011111101100";
        when 5344 => y_in <= "10010100"; x_in <= "01100000"; z_correct<="1101011110000000";
        when 5345 => y_in <= "10010100"; x_in <= "01100001"; z_correct<="1101011100010100";
        when 5346 => y_in <= "10010100"; x_in <= "01100010"; z_correct<="1101011010101000";
        when 5347 => y_in <= "10010100"; x_in <= "01100011"; z_correct<="1101011000111100";
        when 5348 => y_in <= "10010100"; x_in <= "01100100"; z_correct<="1101010111010000";
        when 5349 => y_in <= "10010100"; x_in <= "01100101"; z_correct<="1101010101100100";
        when 5350 => y_in <= "10010100"; x_in <= "01100110"; z_correct<="1101010011111000";
        when 5351 => y_in <= "10010100"; x_in <= "01100111"; z_correct<="1101010010001100";
        when 5352 => y_in <= "10010100"; x_in <= "01101000"; z_correct<="1101010000100000";
        when 5353 => y_in <= "10010100"; x_in <= "01101001"; z_correct<="1101001110110100";
        when 5354 => y_in <= "10010100"; x_in <= "01101010"; z_correct<="1101001101001000";
        when 5355 => y_in <= "10010100"; x_in <= "01101011"; z_correct<="1101001011011100";
        when 5356 => y_in <= "10010100"; x_in <= "01101100"; z_correct<="1101001001110000";
        when 5357 => y_in <= "10010100"; x_in <= "01101101"; z_correct<="1101001000000100";
        when 5358 => y_in <= "10010100"; x_in <= "01101110"; z_correct<="1101000110011000";
        when 5359 => y_in <= "10010100"; x_in <= "01101111"; z_correct<="1101000100101100";
        when 5360 => y_in <= "10010100"; x_in <= "01110000"; z_correct<="1101000011000000";
        when 5361 => y_in <= "10010100"; x_in <= "01110001"; z_correct<="1101000001010100";
        when 5362 => y_in <= "10010100"; x_in <= "01110010"; z_correct<="1100111111101000";
        when 5363 => y_in <= "10010100"; x_in <= "01110011"; z_correct<="1100111101111100";
        when 5364 => y_in <= "10010100"; x_in <= "01110100"; z_correct<="1100111100010000";
        when 5365 => y_in <= "10010100"; x_in <= "01110101"; z_correct<="1100111010100100";
        when 5366 => y_in <= "10010100"; x_in <= "01110110"; z_correct<="1100111000111000";
        when 5367 => y_in <= "10010100"; x_in <= "01110111"; z_correct<="1100110111001100";
        when 5368 => y_in <= "10010100"; x_in <= "01111000"; z_correct<="1100110101100000";
        when 5369 => y_in <= "10010100"; x_in <= "01111001"; z_correct<="1100110011110100";
        when 5370 => y_in <= "10010100"; x_in <= "01111010"; z_correct<="1100110010001000";
        when 5371 => y_in <= "10010100"; x_in <= "01111011"; z_correct<="1100110000011100";
        when 5372 => y_in <= "10010100"; x_in <= "01111100"; z_correct<="1100101110110000";
        when 5373 => y_in <= "10010100"; x_in <= "01111101"; z_correct<="1100101101000100";
        when 5374 => y_in <= "10010100"; x_in <= "01111110"; z_correct<="1100101011011000";
        when 5375 => y_in <= "10010100"; x_in <= "01111111"; z_correct<="1100101001101100";
        when 5376 => y_in <= "10010101"; x_in <= "10000000"; z_correct<="0011010110000000";
        when 5377 => y_in <= "10010101"; x_in <= "10000001"; z_correct<="0011010100010101";
        when 5378 => y_in <= "10010101"; x_in <= "10000010"; z_correct<="0011010010101010";
        when 5379 => y_in <= "10010101"; x_in <= "10000011"; z_correct<="0011010000111111";
        when 5380 => y_in <= "10010101"; x_in <= "10000100"; z_correct<="0011001111010100";
        when 5381 => y_in <= "10010101"; x_in <= "10000101"; z_correct<="0011001101101001";
        when 5382 => y_in <= "10010101"; x_in <= "10000110"; z_correct<="0011001011111110";
        when 5383 => y_in <= "10010101"; x_in <= "10000111"; z_correct<="0011001010010011";
        when 5384 => y_in <= "10010101"; x_in <= "10001000"; z_correct<="0011001000101000";
        when 5385 => y_in <= "10010101"; x_in <= "10001001"; z_correct<="0011000110111101";
        when 5386 => y_in <= "10010101"; x_in <= "10001010"; z_correct<="0011000101010010";
        when 5387 => y_in <= "10010101"; x_in <= "10001011"; z_correct<="0011000011100111";
        when 5388 => y_in <= "10010101"; x_in <= "10001100"; z_correct<="0011000001111100";
        when 5389 => y_in <= "10010101"; x_in <= "10001101"; z_correct<="0011000000010001";
        when 5390 => y_in <= "10010101"; x_in <= "10001110"; z_correct<="0010111110100110";
        when 5391 => y_in <= "10010101"; x_in <= "10001111"; z_correct<="0010111100111011";
        when 5392 => y_in <= "10010101"; x_in <= "10010000"; z_correct<="0010111011010000";
        when 5393 => y_in <= "10010101"; x_in <= "10010001"; z_correct<="0010111001100101";
        when 5394 => y_in <= "10010101"; x_in <= "10010010"; z_correct<="0010110111111010";
        when 5395 => y_in <= "10010101"; x_in <= "10010011"; z_correct<="0010110110001111";
        when 5396 => y_in <= "10010101"; x_in <= "10010100"; z_correct<="0010110100100100";
        when 5397 => y_in <= "10010101"; x_in <= "10010101"; z_correct<="0010110010111001";
        when 5398 => y_in <= "10010101"; x_in <= "10010110"; z_correct<="0010110001001110";
        when 5399 => y_in <= "10010101"; x_in <= "10010111"; z_correct<="0010101111100011";
        when 5400 => y_in <= "10010101"; x_in <= "10011000"; z_correct<="0010101101111000";
        when 5401 => y_in <= "10010101"; x_in <= "10011001"; z_correct<="0010101100001101";
        when 5402 => y_in <= "10010101"; x_in <= "10011010"; z_correct<="0010101010100010";
        when 5403 => y_in <= "10010101"; x_in <= "10011011"; z_correct<="0010101000110111";
        when 5404 => y_in <= "10010101"; x_in <= "10011100"; z_correct<="0010100111001100";
        when 5405 => y_in <= "10010101"; x_in <= "10011101"; z_correct<="0010100101100001";
        when 5406 => y_in <= "10010101"; x_in <= "10011110"; z_correct<="0010100011110110";
        when 5407 => y_in <= "10010101"; x_in <= "10011111"; z_correct<="0010100010001011";
        when 5408 => y_in <= "10010101"; x_in <= "10100000"; z_correct<="0010100000100000";
        when 5409 => y_in <= "10010101"; x_in <= "10100001"; z_correct<="0010011110110101";
        when 5410 => y_in <= "10010101"; x_in <= "10100010"; z_correct<="0010011101001010";
        when 5411 => y_in <= "10010101"; x_in <= "10100011"; z_correct<="0010011011011111";
        when 5412 => y_in <= "10010101"; x_in <= "10100100"; z_correct<="0010011001110100";
        when 5413 => y_in <= "10010101"; x_in <= "10100101"; z_correct<="0010011000001001";
        when 5414 => y_in <= "10010101"; x_in <= "10100110"; z_correct<="0010010110011110";
        when 5415 => y_in <= "10010101"; x_in <= "10100111"; z_correct<="0010010100110011";
        when 5416 => y_in <= "10010101"; x_in <= "10101000"; z_correct<="0010010011001000";
        when 5417 => y_in <= "10010101"; x_in <= "10101001"; z_correct<="0010010001011101";
        when 5418 => y_in <= "10010101"; x_in <= "10101010"; z_correct<="0010001111110010";
        when 5419 => y_in <= "10010101"; x_in <= "10101011"; z_correct<="0010001110000111";
        when 5420 => y_in <= "10010101"; x_in <= "10101100"; z_correct<="0010001100011100";
        when 5421 => y_in <= "10010101"; x_in <= "10101101"; z_correct<="0010001010110001";
        when 5422 => y_in <= "10010101"; x_in <= "10101110"; z_correct<="0010001001000110";
        when 5423 => y_in <= "10010101"; x_in <= "10101111"; z_correct<="0010000111011011";
        when 5424 => y_in <= "10010101"; x_in <= "10110000"; z_correct<="0010000101110000";
        when 5425 => y_in <= "10010101"; x_in <= "10110001"; z_correct<="0010000100000101";
        when 5426 => y_in <= "10010101"; x_in <= "10110010"; z_correct<="0010000010011010";
        when 5427 => y_in <= "10010101"; x_in <= "10110011"; z_correct<="0010000000101111";
        when 5428 => y_in <= "10010101"; x_in <= "10110100"; z_correct<="0001111111000100";
        when 5429 => y_in <= "10010101"; x_in <= "10110101"; z_correct<="0001111101011001";
        when 5430 => y_in <= "10010101"; x_in <= "10110110"; z_correct<="0001111011101110";
        when 5431 => y_in <= "10010101"; x_in <= "10110111"; z_correct<="0001111010000011";
        when 5432 => y_in <= "10010101"; x_in <= "10111000"; z_correct<="0001111000011000";
        when 5433 => y_in <= "10010101"; x_in <= "10111001"; z_correct<="0001110110101101";
        when 5434 => y_in <= "10010101"; x_in <= "10111010"; z_correct<="0001110101000010";
        when 5435 => y_in <= "10010101"; x_in <= "10111011"; z_correct<="0001110011010111";
        when 5436 => y_in <= "10010101"; x_in <= "10111100"; z_correct<="0001110001101100";
        when 5437 => y_in <= "10010101"; x_in <= "10111101"; z_correct<="0001110000000001";
        when 5438 => y_in <= "10010101"; x_in <= "10111110"; z_correct<="0001101110010110";
        when 5439 => y_in <= "10010101"; x_in <= "10111111"; z_correct<="0001101100101011";
        when 5440 => y_in <= "10010101"; x_in <= "11000000"; z_correct<="0001101011000000";
        when 5441 => y_in <= "10010101"; x_in <= "11000001"; z_correct<="0001101001010101";
        when 5442 => y_in <= "10010101"; x_in <= "11000010"; z_correct<="0001100111101010";
        when 5443 => y_in <= "10010101"; x_in <= "11000011"; z_correct<="0001100101111111";
        when 5444 => y_in <= "10010101"; x_in <= "11000100"; z_correct<="0001100100010100";
        when 5445 => y_in <= "10010101"; x_in <= "11000101"; z_correct<="0001100010101001";
        when 5446 => y_in <= "10010101"; x_in <= "11000110"; z_correct<="0001100000111110";
        when 5447 => y_in <= "10010101"; x_in <= "11000111"; z_correct<="0001011111010011";
        when 5448 => y_in <= "10010101"; x_in <= "11001000"; z_correct<="0001011101101000";
        when 5449 => y_in <= "10010101"; x_in <= "11001001"; z_correct<="0001011011111101";
        when 5450 => y_in <= "10010101"; x_in <= "11001010"; z_correct<="0001011010010010";
        when 5451 => y_in <= "10010101"; x_in <= "11001011"; z_correct<="0001011000100111";
        when 5452 => y_in <= "10010101"; x_in <= "11001100"; z_correct<="0001010110111100";
        when 5453 => y_in <= "10010101"; x_in <= "11001101"; z_correct<="0001010101010001";
        when 5454 => y_in <= "10010101"; x_in <= "11001110"; z_correct<="0001010011100110";
        when 5455 => y_in <= "10010101"; x_in <= "11001111"; z_correct<="0001010001111011";
        when 5456 => y_in <= "10010101"; x_in <= "11010000"; z_correct<="0001010000010000";
        when 5457 => y_in <= "10010101"; x_in <= "11010001"; z_correct<="0001001110100101";
        when 5458 => y_in <= "10010101"; x_in <= "11010010"; z_correct<="0001001100111010";
        when 5459 => y_in <= "10010101"; x_in <= "11010011"; z_correct<="0001001011001111";
        when 5460 => y_in <= "10010101"; x_in <= "11010100"; z_correct<="0001001001100100";
        when 5461 => y_in <= "10010101"; x_in <= "11010101"; z_correct<="0001000111111001";
        when 5462 => y_in <= "10010101"; x_in <= "11010110"; z_correct<="0001000110001110";
        when 5463 => y_in <= "10010101"; x_in <= "11010111"; z_correct<="0001000100100011";
        when 5464 => y_in <= "10010101"; x_in <= "11011000"; z_correct<="0001000010111000";
        when 5465 => y_in <= "10010101"; x_in <= "11011001"; z_correct<="0001000001001101";
        when 5466 => y_in <= "10010101"; x_in <= "11011010"; z_correct<="0000111111100010";
        when 5467 => y_in <= "10010101"; x_in <= "11011011"; z_correct<="0000111101110111";
        when 5468 => y_in <= "10010101"; x_in <= "11011100"; z_correct<="0000111100001100";
        when 5469 => y_in <= "10010101"; x_in <= "11011101"; z_correct<="0000111010100001";
        when 5470 => y_in <= "10010101"; x_in <= "11011110"; z_correct<="0000111000110110";
        when 5471 => y_in <= "10010101"; x_in <= "11011111"; z_correct<="0000110111001011";
        when 5472 => y_in <= "10010101"; x_in <= "11100000"; z_correct<="0000110101100000";
        when 5473 => y_in <= "10010101"; x_in <= "11100001"; z_correct<="0000110011110101";
        when 5474 => y_in <= "10010101"; x_in <= "11100010"; z_correct<="0000110010001010";
        when 5475 => y_in <= "10010101"; x_in <= "11100011"; z_correct<="0000110000011111";
        when 5476 => y_in <= "10010101"; x_in <= "11100100"; z_correct<="0000101110110100";
        when 5477 => y_in <= "10010101"; x_in <= "11100101"; z_correct<="0000101101001001";
        when 5478 => y_in <= "10010101"; x_in <= "11100110"; z_correct<="0000101011011110";
        when 5479 => y_in <= "10010101"; x_in <= "11100111"; z_correct<="0000101001110011";
        when 5480 => y_in <= "10010101"; x_in <= "11101000"; z_correct<="0000101000001000";
        when 5481 => y_in <= "10010101"; x_in <= "11101001"; z_correct<="0000100110011101";
        when 5482 => y_in <= "10010101"; x_in <= "11101010"; z_correct<="0000100100110010";
        when 5483 => y_in <= "10010101"; x_in <= "11101011"; z_correct<="0000100011000111";
        when 5484 => y_in <= "10010101"; x_in <= "11101100"; z_correct<="0000100001011100";
        when 5485 => y_in <= "10010101"; x_in <= "11101101"; z_correct<="0000011111110001";
        when 5486 => y_in <= "10010101"; x_in <= "11101110"; z_correct<="0000011110000110";
        when 5487 => y_in <= "10010101"; x_in <= "11101111"; z_correct<="0000011100011011";
        when 5488 => y_in <= "10010101"; x_in <= "11110000"; z_correct<="0000011010110000";
        when 5489 => y_in <= "10010101"; x_in <= "11110001"; z_correct<="0000011001000101";
        when 5490 => y_in <= "10010101"; x_in <= "11110010"; z_correct<="0000010111011010";
        when 5491 => y_in <= "10010101"; x_in <= "11110011"; z_correct<="0000010101101111";
        when 5492 => y_in <= "10010101"; x_in <= "11110100"; z_correct<="0000010100000100";
        when 5493 => y_in <= "10010101"; x_in <= "11110101"; z_correct<="0000010010011001";
        when 5494 => y_in <= "10010101"; x_in <= "11110110"; z_correct<="0000010000101110";
        when 5495 => y_in <= "10010101"; x_in <= "11110111"; z_correct<="0000001111000011";
        when 5496 => y_in <= "10010101"; x_in <= "11111000"; z_correct<="0000001101011000";
        when 5497 => y_in <= "10010101"; x_in <= "11111001"; z_correct<="0000001011101101";
        when 5498 => y_in <= "10010101"; x_in <= "11111010"; z_correct<="0000001010000010";
        when 5499 => y_in <= "10010101"; x_in <= "11111011"; z_correct<="0000001000010111";
        when 5500 => y_in <= "10010101"; x_in <= "11111100"; z_correct<="0000000110101100";
        when 5501 => y_in <= "10010101"; x_in <= "11111101"; z_correct<="0000000101000001";
        when 5502 => y_in <= "10010101"; x_in <= "11111110"; z_correct<="0000000011010110";
        when 5503 => y_in <= "10010101"; x_in <= "11111111"; z_correct<="0000000001101011";
        when 5504 => y_in <= "10010101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 5505 => y_in <= "10010101"; x_in <= "00000001"; z_correct<="1111111110010101";
        when 5506 => y_in <= "10010101"; x_in <= "00000010"; z_correct<="1111111100101010";
        when 5507 => y_in <= "10010101"; x_in <= "00000011"; z_correct<="1111111010111111";
        when 5508 => y_in <= "10010101"; x_in <= "00000100"; z_correct<="1111111001010100";
        when 5509 => y_in <= "10010101"; x_in <= "00000101"; z_correct<="1111110111101001";
        when 5510 => y_in <= "10010101"; x_in <= "00000110"; z_correct<="1111110101111110";
        when 5511 => y_in <= "10010101"; x_in <= "00000111"; z_correct<="1111110100010011";
        when 5512 => y_in <= "10010101"; x_in <= "00001000"; z_correct<="1111110010101000";
        when 5513 => y_in <= "10010101"; x_in <= "00001001"; z_correct<="1111110000111101";
        when 5514 => y_in <= "10010101"; x_in <= "00001010"; z_correct<="1111101111010010";
        when 5515 => y_in <= "10010101"; x_in <= "00001011"; z_correct<="1111101101100111";
        when 5516 => y_in <= "10010101"; x_in <= "00001100"; z_correct<="1111101011111100";
        when 5517 => y_in <= "10010101"; x_in <= "00001101"; z_correct<="1111101010010001";
        when 5518 => y_in <= "10010101"; x_in <= "00001110"; z_correct<="1111101000100110";
        when 5519 => y_in <= "10010101"; x_in <= "00001111"; z_correct<="1111100110111011";
        when 5520 => y_in <= "10010101"; x_in <= "00010000"; z_correct<="1111100101010000";
        when 5521 => y_in <= "10010101"; x_in <= "00010001"; z_correct<="1111100011100101";
        when 5522 => y_in <= "10010101"; x_in <= "00010010"; z_correct<="1111100001111010";
        when 5523 => y_in <= "10010101"; x_in <= "00010011"; z_correct<="1111100000001111";
        when 5524 => y_in <= "10010101"; x_in <= "00010100"; z_correct<="1111011110100100";
        when 5525 => y_in <= "10010101"; x_in <= "00010101"; z_correct<="1111011100111001";
        when 5526 => y_in <= "10010101"; x_in <= "00010110"; z_correct<="1111011011001110";
        when 5527 => y_in <= "10010101"; x_in <= "00010111"; z_correct<="1111011001100011";
        when 5528 => y_in <= "10010101"; x_in <= "00011000"; z_correct<="1111010111111000";
        when 5529 => y_in <= "10010101"; x_in <= "00011001"; z_correct<="1111010110001101";
        when 5530 => y_in <= "10010101"; x_in <= "00011010"; z_correct<="1111010100100010";
        when 5531 => y_in <= "10010101"; x_in <= "00011011"; z_correct<="1111010010110111";
        when 5532 => y_in <= "10010101"; x_in <= "00011100"; z_correct<="1111010001001100";
        when 5533 => y_in <= "10010101"; x_in <= "00011101"; z_correct<="1111001111100001";
        when 5534 => y_in <= "10010101"; x_in <= "00011110"; z_correct<="1111001101110110";
        when 5535 => y_in <= "10010101"; x_in <= "00011111"; z_correct<="1111001100001011";
        when 5536 => y_in <= "10010101"; x_in <= "00100000"; z_correct<="1111001010100000";
        when 5537 => y_in <= "10010101"; x_in <= "00100001"; z_correct<="1111001000110101";
        when 5538 => y_in <= "10010101"; x_in <= "00100010"; z_correct<="1111000111001010";
        when 5539 => y_in <= "10010101"; x_in <= "00100011"; z_correct<="1111000101011111";
        when 5540 => y_in <= "10010101"; x_in <= "00100100"; z_correct<="1111000011110100";
        when 5541 => y_in <= "10010101"; x_in <= "00100101"; z_correct<="1111000010001001";
        when 5542 => y_in <= "10010101"; x_in <= "00100110"; z_correct<="1111000000011110";
        when 5543 => y_in <= "10010101"; x_in <= "00100111"; z_correct<="1110111110110011";
        when 5544 => y_in <= "10010101"; x_in <= "00101000"; z_correct<="1110111101001000";
        when 5545 => y_in <= "10010101"; x_in <= "00101001"; z_correct<="1110111011011101";
        when 5546 => y_in <= "10010101"; x_in <= "00101010"; z_correct<="1110111001110010";
        when 5547 => y_in <= "10010101"; x_in <= "00101011"; z_correct<="1110111000000111";
        when 5548 => y_in <= "10010101"; x_in <= "00101100"; z_correct<="1110110110011100";
        when 5549 => y_in <= "10010101"; x_in <= "00101101"; z_correct<="1110110100110001";
        when 5550 => y_in <= "10010101"; x_in <= "00101110"; z_correct<="1110110011000110";
        when 5551 => y_in <= "10010101"; x_in <= "00101111"; z_correct<="1110110001011011";
        when 5552 => y_in <= "10010101"; x_in <= "00110000"; z_correct<="1110101111110000";
        when 5553 => y_in <= "10010101"; x_in <= "00110001"; z_correct<="1110101110000101";
        when 5554 => y_in <= "10010101"; x_in <= "00110010"; z_correct<="1110101100011010";
        when 5555 => y_in <= "10010101"; x_in <= "00110011"; z_correct<="1110101010101111";
        when 5556 => y_in <= "10010101"; x_in <= "00110100"; z_correct<="1110101001000100";
        when 5557 => y_in <= "10010101"; x_in <= "00110101"; z_correct<="1110100111011001";
        when 5558 => y_in <= "10010101"; x_in <= "00110110"; z_correct<="1110100101101110";
        when 5559 => y_in <= "10010101"; x_in <= "00110111"; z_correct<="1110100100000011";
        when 5560 => y_in <= "10010101"; x_in <= "00111000"; z_correct<="1110100010011000";
        when 5561 => y_in <= "10010101"; x_in <= "00111001"; z_correct<="1110100000101101";
        when 5562 => y_in <= "10010101"; x_in <= "00111010"; z_correct<="1110011111000010";
        when 5563 => y_in <= "10010101"; x_in <= "00111011"; z_correct<="1110011101010111";
        when 5564 => y_in <= "10010101"; x_in <= "00111100"; z_correct<="1110011011101100";
        when 5565 => y_in <= "10010101"; x_in <= "00111101"; z_correct<="1110011010000001";
        when 5566 => y_in <= "10010101"; x_in <= "00111110"; z_correct<="1110011000010110";
        when 5567 => y_in <= "10010101"; x_in <= "00111111"; z_correct<="1110010110101011";
        when 5568 => y_in <= "10010101"; x_in <= "01000000"; z_correct<="1110010101000000";
        when 5569 => y_in <= "10010101"; x_in <= "01000001"; z_correct<="1110010011010101";
        when 5570 => y_in <= "10010101"; x_in <= "01000010"; z_correct<="1110010001101010";
        when 5571 => y_in <= "10010101"; x_in <= "01000011"; z_correct<="1110001111111111";
        when 5572 => y_in <= "10010101"; x_in <= "01000100"; z_correct<="1110001110010100";
        when 5573 => y_in <= "10010101"; x_in <= "01000101"; z_correct<="1110001100101001";
        when 5574 => y_in <= "10010101"; x_in <= "01000110"; z_correct<="1110001010111110";
        when 5575 => y_in <= "10010101"; x_in <= "01000111"; z_correct<="1110001001010011";
        when 5576 => y_in <= "10010101"; x_in <= "01001000"; z_correct<="1110000111101000";
        when 5577 => y_in <= "10010101"; x_in <= "01001001"; z_correct<="1110000101111101";
        when 5578 => y_in <= "10010101"; x_in <= "01001010"; z_correct<="1110000100010010";
        when 5579 => y_in <= "10010101"; x_in <= "01001011"; z_correct<="1110000010100111";
        when 5580 => y_in <= "10010101"; x_in <= "01001100"; z_correct<="1110000000111100";
        when 5581 => y_in <= "10010101"; x_in <= "01001101"; z_correct<="1101111111010001";
        when 5582 => y_in <= "10010101"; x_in <= "01001110"; z_correct<="1101111101100110";
        when 5583 => y_in <= "10010101"; x_in <= "01001111"; z_correct<="1101111011111011";
        when 5584 => y_in <= "10010101"; x_in <= "01010000"; z_correct<="1101111010010000";
        when 5585 => y_in <= "10010101"; x_in <= "01010001"; z_correct<="1101111000100101";
        when 5586 => y_in <= "10010101"; x_in <= "01010010"; z_correct<="1101110110111010";
        when 5587 => y_in <= "10010101"; x_in <= "01010011"; z_correct<="1101110101001111";
        when 5588 => y_in <= "10010101"; x_in <= "01010100"; z_correct<="1101110011100100";
        when 5589 => y_in <= "10010101"; x_in <= "01010101"; z_correct<="1101110001111001";
        when 5590 => y_in <= "10010101"; x_in <= "01010110"; z_correct<="1101110000001110";
        when 5591 => y_in <= "10010101"; x_in <= "01010111"; z_correct<="1101101110100011";
        when 5592 => y_in <= "10010101"; x_in <= "01011000"; z_correct<="1101101100111000";
        when 5593 => y_in <= "10010101"; x_in <= "01011001"; z_correct<="1101101011001101";
        when 5594 => y_in <= "10010101"; x_in <= "01011010"; z_correct<="1101101001100010";
        when 5595 => y_in <= "10010101"; x_in <= "01011011"; z_correct<="1101100111110111";
        when 5596 => y_in <= "10010101"; x_in <= "01011100"; z_correct<="1101100110001100";
        when 5597 => y_in <= "10010101"; x_in <= "01011101"; z_correct<="1101100100100001";
        when 5598 => y_in <= "10010101"; x_in <= "01011110"; z_correct<="1101100010110110";
        when 5599 => y_in <= "10010101"; x_in <= "01011111"; z_correct<="1101100001001011";
        when 5600 => y_in <= "10010101"; x_in <= "01100000"; z_correct<="1101011111100000";
        when 5601 => y_in <= "10010101"; x_in <= "01100001"; z_correct<="1101011101110101";
        when 5602 => y_in <= "10010101"; x_in <= "01100010"; z_correct<="1101011100001010";
        when 5603 => y_in <= "10010101"; x_in <= "01100011"; z_correct<="1101011010011111";
        when 5604 => y_in <= "10010101"; x_in <= "01100100"; z_correct<="1101011000110100";
        when 5605 => y_in <= "10010101"; x_in <= "01100101"; z_correct<="1101010111001001";
        when 5606 => y_in <= "10010101"; x_in <= "01100110"; z_correct<="1101010101011110";
        when 5607 => y_in <= "10010101"; x_in <= "01100111"; z_correct<="1101010011110011";
        when 5608 => y_in <= "10010101"; x_in <= "01101000"; z_correct<="1101010010001000";
        when 5609 => y_in <= "10010101"; x_in <= "01101001"; z_correct<="1101010000011101";
        when 5610 => y_in <= "10010101"; x_in <= "01101010"; z_correct<="1101001110110010";
        when 5611 => y_in <= "10010101"; x_in <= "01101011"; z_correct<="1101001101000111";
        when 5612 => y_in <= "10010101"; x_in <= "01101100"; z_correct<="1101001011011100";
        when 5613 => y_in <= "10010101"; x_in <= "01101101"; z_correct<="1101001001110001";
        when 5614 => y_in <= "10010101"; x_in <= "01101110"; z_correct<="1101001000000110";
        when 5615 => y_in <= "10010101"; x_in <= "01101111"; z_correct<="1101000110011011";
        when 5616 => y_in <= "10010101"; x_in <= "01110000"; z_correct<="1101000100110000";
        when 5617 => y_in <= "10010101"; x_in <= "01110001"; z_correct<="1101000011000101";
        when 5618 => y_in <= "10010101"; x_in <= "01110010"; z_correct<="1101000001011010";
        when 5619 => y_in <= "10010101"; x_in <= "01110011"; z_correct<="1100111111101111";
        when 5620 => y_in <= "10010101"; x_in <= "01110100"; z_correct<="1100111110000100";
        when 5621 => y_in <= "10010101"; x_in <= "01110101"; z_correct<="1100111100011001";
        when 5622 => y_in <= "10010101"; x_in <= "01110110"; z_correct<="1100111010101110";
        when 5623 => y_in <= "10010101"; x_in <= "01110111"; z_correct<="1100111001000011";
        when 5624 => y_in <= "10010101"; x_in <= "01111000"; z_correct<="1100110111011000";
        when 5625 => y_in <= "10010101"; x_in <= "01111001"; z_correct<="1100110101101101";
        when 5626 => y_in <= "10010101"; x_in <= "01111010"; z_correct<="1100110100000010";
        when 5627 => y_in <= "10010101"; x_in <= "01111011"; z_correct<="1100110010010111";
        when 5628 => y_in <= "10010101"; x_in <= "01111100"; z_correct<="1100110000101100";
        when 5629 => y_in <= "10010101"; x_in <= "01111101"; z_correct<="1100101111000001";
        when 5630 => y_in <= "10010101"; x_in <= "01111110"; z_correct<="1100101101010110";
        when 5631 => y_in <= "10010101"; x_in <= "01111111"; z_correct<="1100101011101011";
        when 5632 => y_in <= "10010110"; x_in <= "10000000"; z_correct<="0011010100000000";
        when 5633 => y_in <= "10010110"; x_in <= "10000001"; z_correct<="0011010010010110";
        when 5634 => y_in <= "10010110"; x_in <= "10000010"; z_correct<="0011010000101100";
        when 5635 => y_in <= "10010110"; x_in <= "10000011"; z_correct<="0011001111000010";
        when 5636 => y_in <= "10010110"; x_in <= "10000100"; z_correct<="0011001101011000";
        when 5637 => y_in <= "10010110"; x_in <= "10000101"; z_correct<="0011001011101110";
        when 5638 => y_in <= "10010110"; x_in <= "10000110"; z_correct<="0011001010000100";
        when 5639 => y_in <= "10010110"; x_in <= "10000111"; z_correct<="0011001000011010";
        when 5640 => y_in <= "10010110"; x_in <= "10001000"; z_correct<="0011000110110000";
        when 5641 => y_in <= "10010110"; x_in <= "10001001"; z_correct<="0011000101000110";
        when 5642 => y_in <= "10010110"; x_in <= "10001010"; z_correct<="0011000011011100";
        when 5643 => y_in <= "10010110"; x_in <= "10001011"; z_correct<="0011000001110010";
        when 5644 => y_in <= "10010110"; x_in <= "10001100"; z_correct<="0011000000001000";
        when 5645 => y_in <= "10010110"; x_in <= "10001101"; z_correct<="0010111110011110";
        when 5646 => y_in <= "10010110"; x_in <= "10001110"; z_correct<="0010111100110100";
        when 5647 => y_in <= "10010110"; x_in <= "10001111"; z_correct<="0010111011001010";
        when 5648 => y_in <= "10010110"; x_in <= "10010000"; z_correct<="0010111001100000";
        when 5649 => y_in <= "10010110"; x_in <= "10010001"; z_correct<="0010110111110110";
        when 5650 => y_in <= "10010110"; x_in <= "10010010"; z_correct<="0010110110001100";
        when 5651 => y_in <= "10010110"; x_in <= "10010011"; z_correct<="0010110100100010";
        when 5652 => y_in <= "10010110"; x_in <= "10010100"; z_correct<="0010110010111000";
        when 5653 => y_in <= "10010110"; x_in <= "10010101"; z_correct<="0010110001001110";
        when 5654 => y_in <= "10010110"; x_in <= "10010110"; z_correct<="0010101111100100";
        when 5655 => y_in <= "10010110"; x_in <= "10010111"; z_correct<="0010101101111010";
        when 5656 => y_in <= "10010110"; x_in <= "10011000"; z_correct<="0010101100010000";
        when 5657 => y_in <= "10010110"; x_in <= "10011001"; z_correct<="0010101010100110";
        when 5658 => y_in <= "10010110"; x_in <= "10011010"; z_correct<="0010101000111100";
        when 5659 => y_in <= "10010110"; x_in <= "10011011"; z_correct<="0010100111010010";
        when 5660 => y_in <= "10010110"; x_in <= "10011100"; z_correct<="0010100101101000";
        when 5661 => y_in <= "10010110"; x_in <= "10011101"; z_correct<="0010100011111110";
        when 5662 => y_in <= "10010110"; x_in <= "10011110"; z_correct<="0010100010010100";
        when 5663 => y_in <= "10010110"; x_in <= "10011111"; z_correct<="0010100000101010";
        when 5664 => y_in <= "10010110"; x_in <= "10100000"; z_correct<="0010011111000000";
        when 5665 => y_in <= "10010110"; x_in <= "10100001"; z_correct<="0010011101010110";
        when 5666 => y_in <= "10010110"; x_in <= "10100010"; z_correct<="0010011011101100";
        when 5667 => y_in <= "10010110"; x_in <= "10100011"; z_correct<="0010011010000010";
        when 5668 => y_in <= "10010110"; x_in <= "10100100"; z_correct<="0010011000011000";
        when 5669 => y_in <= "10010110"; x_in <= "10100101"; z_correct<="0010010110101110";
        when 5670 => y_in <= "10010110"; x_in <= "10100110"; z_correct<="0010010101000100";
        when 5671 => y_in <= "10010110"; x_in <= "10100111"; z_correct<="0010010011011010";
        when 5672 => y_in <= "10010110"; x_in <= "10101000"; z_correct<="0010010001110000";
        when 5673 => y_in <= "10010110"; x_in <= "10101001"; z_correct<="0010010000000110";
        when 5674 => y_in <= "10010110"; x_in <= "10101010"; z_correct<="0010001110011100";
        when 5675 => y_in <= "10010110"; x_in <= "10101011"; z_correct<="0010001100110010";
        when 5676 => y_in <= "10010110"; x_in <= "10101100"; z_correct<="0010001011001000";
        when 5677 => y_in <= "10010110"; x_in <= "10101101"; z_correct<="0010001001011110";
        when 5678 => y_in <= "10010110"; x_in <= "10101110"; z_correct<="0010000111110100";
        when 5679 => y_in <= "10010110"; x_in <= "10101111"; z_correct<="0010000110001010";
        when 5680 => y_in <= "10010110"; x_in <= "10110000"; z_correct<="0010000100100000";
        when 5681 => y_in <= "10010110"; x_in <= "10110001"; z_correct<="0010000010110110";
        when 5682 => y_in <= "10010110"; x_in <= "10110010"; z_correct<="0010000001001100";
        when 5683 => y_in <= "10010110"; x_in <= "10110011"; z_correct<="0001111111100010";
        when 5684 => y_in <= "10010110"; x_in <= "10110100"; z_correct<="0001111101111000";
        when 5685 => y_in <= "10010110"; x_in <= "10110101"; z_correct<="0001111100001110";
        when 5686 => y_in <= "10010110"; x_in <= "10110110"; z_correct<="0001111010100100";
        when 5687 => y_in <= "10010110"; x_in <= "10110111"; z_correct<="0001111000111010";
        when 5688 => y_in <= "10010110"; x_in <= "10111000"; z_correct<="0001110111010000";
        when 5689 => y_in <= "10010110"; x_in <= "10111001"; z_correct<="0001110101100110";
        when 5690 => y_in <= "10010110"; x_in <= "10111010"; z_correct<="0001110011111100";
        when 5691 => y_in <= "10010110"; x_in <= "10111011"; z_correct<="0001110010010010";
        when 5692 => y_in <= "10010110"; x_in <= "10111100"; z_correct<="0001110000101000";
        when 5693 => y_in <= "10010110"; x_in <= "10111101"; z_correct<="0001101110111110";
        when 5694 => y_in <= "10010110"; x_in <= "10111110"; z_correct<="0001101101010100";
        when 5695 => y_in <= "10010110"; x_in <= "10111111"; z_correct<="0001101011101010";
        when 5696 => y_in <= "10010110"; x_in <= "11000000"; z_correct<="0001101010000000";
        when 5697 => y_in <= "10010110"; x_in <= "11000001"; z_correct<="0001101000010110";
        when 5698 => y_in <= "10010110"; x_in <= "11000010"; z_correct<="0001100110101100";
        when 5699 => y_in <= "10010110"; x_in <= "11000011"; z_correct<="0001100101000010";
        when 5700 => y_in <= "10010110"; x_in <= "11000100"; z_correct<="0001100011011000";
        when 5701 => y_in <= "10010110"; x_in <= "11000101"; z_correct<="0001100001101110";
        when 5702 => y_in <= "10010110"; x_in <= "11000110"; z_correct<="0001100000000100";
        when 5703 => y_in <= "10010110"; x_in <= "11000111"; z_correct<="0001011110011010";
        when 5704 => y_in <= "10010110"; x_in <= "11001000"; z_correct<="0001011100110000";
        when 5705 => y_in <= "10010110"; x_in <= "11001001"; z_correct<="0001011011000110";
        when 5706 => y_in <= "10010110"; x_in <= "11001010"; z_correct<="0001011001011100";
        when 5707 => y_in <= "10010110"; x_in <= "11001011"; z_correct<="0001010111110010";
        when 5708 => y_in <= "10010110"; x_in <= "11001100"; z_correct<="0001010110001000";
        when 5709 => y_in <= "10010110"; x_in <= "11001101"; z_correct<="0001010100011110";
        when 5710 => y_in <= "10010110"; x_in <= "11001110"; z_correct<="0001010010110100";
        when 5711 => y_in <= "10010110"; x_in <= "11001111"; z_correct<="0001010001001010";
        when 5712 => y_in <= "10010110"; x_in <= "11010000"; z_correct<="0001001111100000";
        when 5713 => y_in <= "10010110"; x_in <= "11010001"; z_correct<="0001001101110110";
        when 5714 => y_in <= "10010110"; x_in <= "11010010"; z_correct<="0001001100001100";
        when 5715 => y_in <= "10010110"; x_in <= "11010011"; z_correct<="0001001010100010";
        when 5716 => y_in <= "10010110"; x_in <= "11010100"; z_correct<="0001001000111000";
        when 5717 => y_in <= "10010110"; x_in <= "11010101"; z_correct<="0001000111001110";
        when 5718 => y_in <= "10010110"; x_in <= "11010110"; z_correct<="0001000101100100";
        when 5719 => y_in <= "10010110"; x_in <= "11010111"; z_correct<="0001000011111010";
        when 5720 => y_in <= "10010110"; x_in <= "11011000"; z_correct<="0001000010010000";
        when 5721 => y_in <= "10010110"; x_in <= "11011001"; z_correct<="0001000000100110";
        when 5722 => y_in <= "10010110"; x_in <= "11011010"; z_correct<="0000111110111100";
        when 5723 => y_in <= "10010110"; x_in <= "11011011"; z_correct<="0000111101010010";
        when 5724 => y_in <= "10010110"; x_in <= "11011100"; z_correct<="0000111011101000";
        when 5725 => y_in <= "10010110"; x_in <= "11011101"; z_correct<="0000111001111110";
        when 5726 => y_in <= "10010110"; x_in <= "11011110"; z_correct<="0000111000010100";
        when 5727 => y_in <= "10010110"; x_in <= "11011111"; z_correct<="0000110110101010";
        when 5728 => y_in <= "10010110"; x_in <= "11100000"; z_correct<="0000110101000000";
        when 5729 => y_in <= "10010110"; x_in <= "11100001"; z_correct<="0000110011010110";
        when 5730 => y_in <= "10010110"; x_in <= "11100010"; z_correct<="0000110001101100";
        when 5731 => y_in <= "10010110"; x_in <= "11100011"; z_correct<="0000110000000010";
        when 5732 => y_in <= "10010110"; x_in <= "11100100"; z_correct<="0000101110011000";
        when 5733 => y_in <= "10010110"; x_in <= "11100101"; z_correct<="0000101100101110";
        when 5734 => y_in <= "10010110"; x_in <= "11100110"; z_correct<="0000101011000100";
        when 5735 => y_in <= "10010110"; x_in <= "11100111"; z_correct<="0000101001011010";
        when 5736 => y_in <= "10010110"; x_in <= "11101000"; z_correct<="0000100111110000";
        when 5737 => y_in <= "10010110"; x_in <= "11101001"; z_correct<="0000100110000110";
        when 5738 => y_in <= "10010110"; x_in <= "11101010"; z_correct<="0000100100011100";
        when 5739 => y_in <= "10010110"; x_in <= "11101011"; z_correct<="0000100010110010";
        when 5740 => y_in <= "10010110"; x_in <= "11101100"; z_correct<="0000100001001000";
        when 5741 => y_in <= "10010110"; x_in <= "11101101"; z_correct<="0000011111011110";
        when 5742 => y_in <= "10010110"; x_in <= "11101110"; z_correct<="0000011101110100";
        when 5743 => y_in <= "10010110"; x_in <= "11101111"; z_correct<="0000011100001010";
        when 5744 => y_in <= "10010110"; x_in <= "11110000"; z_correct<="0000011010100000";
        when 5745 => y_in <= "10010110"; x_in <= "11110001"; z_correct<="0000011000110110";
        when 5746 => y_in <= "10010110"; x_in <= "11110010"; z_correct<="0000010111001100";
        when 5747 => y_in <= "10010110"; x_in <= "11110011"; z_correct<="0000010101100010";
        when 5748 => y_in <= "10010110"; x_in <= "11110100"; z_correct<="0000010011111000";
        when 5749 => y_in <= "10010110"; x_in <= "11110101"; z_correct<="0000010010001110";
        when 5750 => y_in <= "10010110"; x_in <= "11110110"; z_correct<="0000010000100100";
        when 5751 => y_in <= "10010110"; x_in <= "11110111"; z_correct<="0000001110111010";
        when 5752 => y_in <= "10010110"; x_in <= "11111000"; z_correct<="0000001101010000";
        when 5753 => y_in <= "10010110"; x_in <= "11111001"; z_correct<="0000001011100110";
        when 5754 => y_in <= "10010110"; x_in <= "11111010"; z_correct<="0000001001111100";
        when 5755 => y_in <= "10010110"; x_in <= "11111011"; z_correct<="0000001000010010";
        when 5756 => y_in <= "10010110"; x_in <= "11111100"; z_correct<="0000000110101000";
        when 5757 => y_in <= "10010110"; x_in <= "11111101"; z_correct<="0000000100111110";
        when 5758 => y_in <= "10010110"; x_in <= "11111110"; z_correct<="0000000011010100";
        when 5759 => y_in <= "10010110"; x_in <= "11111111"; z_correct<="0000000001101010";
        when 5760 => y_in <= "10010110"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 5761 => y_in <= "10010110"; x_in <= "00000001"; z_correct<="1111111110010110";
        when 5762 => y_in <= "10010110"; x_in <= "00000010"; z_correct<="1111111100101100";
        when 5763 => y_in <= "10010110"; x_in <= "00000011"; z_correct<="1111111011000010";
        when 5764 => y_in <= "10010110"; x_in <= "00000100"; z_correct<="1111111001011000";
        when 5765 => y_in <= "10010110"; x_in <= "00000101"; z_correct<="1111110111101110";
        when 5766 => y_in <= "10010110"; x_in <= "00000110"; z_correct<="1111110110000100";
        when 5767 => y_in <= "10010110"; x_in <= "00000111"; z_correct<="1111110100011010";
        when 5768 => y_in <= "10010110"; x_in <= "00001000"; z_correct<="1111110010110000";
        when 5769 => y_in <= "10010110"; x_in <= "00001001"; z_correct<="1111110001000110";
        when 5770 => y_in <= "10010110"; x_in <= "00001010"; z_correct<="1111101111011100";
        when 5771 => y_in <= "10010110"; x_in <= "00001011"; z_correct<="1111101101110010";
        when 5772 => y_in <= "10010110"; x_in <= "00001100"; z_correct<="1111101100001000";
        when 5773 => y_in <= "10010110"; x_in <= "00001101"; z_correct<="1111101010011110";
        when 5774 => y_in <= "10010110"; x_in <= "00001110"; z_correct<="1111101000110100";
        when 5775 => y_in <= "10010110"; x_in <= "00001111"; z_correct<="1111100111001010";
        when 5776 => y_in <= "10010110"; x_in <= "00010000"; z_correct<="1111100101100000";
        when 5777 => y_in <= "10010110"; x_in <= "00010001"; z_correct<="1111100011110110";
        when 5778 => y_in <= "10010110"; x_in <= "00010010"; z_correct<="1111100010001100";
        when 5779 => y_in <= "10010110"; x_in <= "00010011"; z_correct<="1111100000100010";
        when 5780 => y_in <= "10010110"; x_in <= "00010100"; z_correct<="1111011110111000";
        when 5781 => y_in <= "10010110"; x_in <= "00010101"; z_correct<="1111011101001110";
        when 5782 => y_in <= "10010110"; x_in <= "00010110"; z_correct<="1111011011100100";
        when 5783 => y_in <= "10010110"; x_in <= "00010111"; z_correct<="1111011001111010";
        when 5784 => y_in <= "10010110"; x_in <= "00011000"; z_correct<="1111011000010000";
        when 5785 => y_in <= "10010110"; x_in <= "00011001"; z_correct<="1111010110100110";
        when 5786 => y_in <= "10010110"; x_in <= "00011010"; z_correct<="1111010100111100";
        when 5787 => y_in <= "10010110"; x_in <= "00011011"; z_correct<="1111010011010010";
        when 5788 => y_in <= "10010110"; x_in <= "00011100"; z_correct<="1111010001101000";
        when 5789 => y_in <= "10010110"; x_in <= "00011101"; z_correct<="1111001111111110";
        when 5790 => y_in <= "10010110"; x_in <= "00011110"; z_correct<="1111001110010100";
        when 5791 => y_in <= "10010110"; x_in <= "00011111"; z_correct<="1111001100101010";
        when 5792 => y_in <= "10010110"; x_in <= "00100000"; z_correct<="1111001011000000";
        when 5793 => y_in <= "10010110"; x_in <= "00100001"; z_correct<="1111001001010110";
        when 5794 => y_in <= "10010110"; x_in <= "00100010"; z_correct<="1111000111101100";
        when 5795 => y_in <= "10010110"; x_in <= "00100011"; z_correct<="1111000110000010";
        when 5796 => y_in <= "10010110"; x_in <= "00100100"; z_correct<="1111000100011000";
        when 5797 => y_in <= "10010110"; x_in <= "00100101"; z_correct<="1111000010101110";
        when 5798 => y_in <= "10010110"; x_in <= "00100110"; z_correct<="1111000001000100";
        when 5799 => y_in <= "10010110"; x_in <= "00100111"; z_correct<="1110111111011010";
        when 5800 => y_in <= "10010110"; x_in <= "00101000"; z_correct<="1110111101110000";
        when 5801 => y_in <= "10010110"; x_in <= "00101001"; z_correct<="1110111100000110";
        when 5802 => y_in <= "10010110"; x_in <= "00101010"; z_correct<="1110111010011100";
        when 5803 => y_in <= "10010110"; x_in <= "00101011"; z_correct<="1110111000110010";
        when 5804 => y_in <= "10010110"; x_in <= "00101100"; z_correct<="1110110111001000";
        when 5805 => y_in <= "10010110"; x_in <= "00101101"; z_correct<="1110110101011110";
        when 5806 => y_in <= "10010110"; x_in <= "00101110"; z_correct<="1110110011110100";
        when 5807 => y_in <= "10010110"; x_in <= "00101111"; z_correct<="1110110010001010";
        when 5808 => y_in <= "10010110"; x_in <= "00110000"; z_correct<="1110110000100000";
        when 5809 => y_in <= "10010110"; x_in <= "00110001"; z_correct<="1110101110110110";
        when 5810 => y_in <= "10010110"; x_in <= "00110010"; z_correct<="1110101101001100";
        when 5811 => y_in <= "10010110"; x_in <= "00110011"; z_correct<="1110101011100010";
        when 5812 => y_in <= "10010110"; x_in <= "00110100"; z_correct<="1110101001111000";
        when 5813 => y_in <= "10010110"; x_in <= "00110101"; z_correct<="1110101000001110";
        when 5814 => y_in <= "10010110"; x_in <= "00110110"; z_correct<="1110100110100100";
        when 5815 => y_in <= "10010110"; x_in <= "00110111"; z_correct<="1110100100111010";
        when 5816 => y_in <= "10010110"; x_in <= "00111000"; z_correct<="1110100011010000";
        when 5817 => y_in <= "10010110"; x_in <= "00111001"; z_correct<="1110100001100110";
        when 5818 => y_in <= "10010110"; x_in <= "00111010"; z_correct<="1110011111111100";
        when 5819 => y_in <= "10010110"; x_in <= "00111011"; z_correct<="1110011110010010";
        when 5820 => y_in <= "10010110"; x_in <= "00111100"; z_correct<="1110011100101000";
        when 5821 => y_in <= "10010110"; x_in <= "00111101"; z_correct<="1110011010111110";
        when 5822 => y_in <= "10010110"; x_in <= "00111110"; z_correct<="1110011001010100";
        when 5823 => y_in <= "10010110"; x_in <= "00111111"; z_correct<="1110010111101010";
        when 5824 => y_in <= "10010110"; x_in <= "01000000"; z_correct<="1110010110000000";
        when 5825 => y_in <= "10010110"; x_in <= "01000001"; z_correct<="1110010100010110";
        when 5826 => y_in <= "10010110"; x_in <= "01000010"; z_correct<="1110010010101100";
        when 5827 => y_in <= "10010110"; x_in <= "01000011"; z_correct<="1110010001000010";
        when 5828 => y_in <= "10010110"; x_in <= "01000100"; z_correct<="1110001111011000";
        when 5829 => y_in <= "10010110"; x_in <= "01000101"; z_correct<="1110001101101110";
        when 5830 => y_in <= "10010110"; x_in <= "01000110"; z_correct<="1110001100000100";
        when 5831 => y_in <= "10010110"; x_in <= "01000111"; z_correct<="1110001010011010";
        when 5832 => y_in <= "10010110"; x_in <= "01001000"; z_correct<="1110001000110000";
        when 5833 => y_in <= "10010110"; x_in <= "01001001"; z_correct<="1110000111000110";
        when 5834 => y_in <= "10010110"; x_in <= "01001010"; z_correct<="1110000101011100";
        when 5835 => y_in <= "10010110"; x_in <= "01001011"; z_correct<="1110000011110010";
        when 5836 => y_in <= "10010110"; x_in <= "01001100"; z_correct<="1110000010001000";
        when 5837 => y_in <= "10010110"; x_in <= "01001101"; z_correct<="1110000000011110";
        when 5838 => y_in <= "10010110"; x_in <= "01001110"; z_correct<="1101111110110100";
        when 5839 => y_in <= "10010110"; x_in <= "01001111"; z_correct<="1101111101001010";
        when 5840 => y_in <= "10010110"; x_in <= "01010000"; z_correct<="1101111011100000";
        when 5841 => y_in <= "10010110"; x_in <= "01010001"; z_correct<="1101111001110110";
        when 5842 => y_in <= "10010110"; x_in <= "01010010"; z_correct<="1101111000001100";
        when 5843 => y_in <= "10010110"; x_in <= "01010011"; z_correct<="1101110110100010";
        when 5844 => y_in <= "10010110"; x_in <= "01010100"; z_correct<="1101110100111000";
        when 5845 => y_in <= "10010110"; x_in <= "01010101"; z_correct<="1101110011001110";
        when 5846 => y_in <= "10010110"; x_in <= "01010110"; z_correct<="1101110001100100";
        when 5847 => y_in <= "10010110"; x_in <= "01010111"; z_correct<="1101101111111010";
        when 5848 => y_in <= "10010110"; x_in <= "01011000"; z_correct<="1101101110010000";
        when 5849 => y_in <= "10010110"; x_in <= "01011001"; z_correct<="1101101100100110";
        when 5850 => y_in <= "10010110"; x_in <= "01011010"; z_correct<="1101101010111100";
        when 5851 => y_in <= "10010110"; x_in <= "01011011"; z_correct<="1101101001010010";
        when 5852 => y_in <= "10010110"; x_in <= "01011100"; z_correct<="1101100111101000";
        when 5853 => y_in <= "10010110"; x_in <= "01011101"; z_correct<="1101100101111110";
        when 5854 => y_in <= "10010110"; x_in <= "01011110"; z_correct<="1101100100010100";
        when 5855 => y_in <= "10010110"; x_in <= "01011111"; z_correct<="1101100010101010";
        when 5856 => y_in <= "10010110"; x_in <= "01100000"; z_correct<="1101100001000000";
        when 5857 => y_in <= "10010110"; x_in <= "01100001"; z_correct<="1101011111010110";
        when 5858 => y_in <= "10010110"; x_in <= "01100010"; z_correct<="1101011101101100";
        when 5859 => y_in <= "10010110"; x_in <= "01100011"; z_correct<="1101011100000010";
        when 5860 => y_in <= "10010110"; x_in <= "01100100"; z_correct<="1101011010011000";
        when 5861 => y_in <= "10010110"; x_in <= "01100101"; z_correct<="1101011000101110";
        when 5862 => y_in <= "10010110"; x_in <= "01100110"; z_correct<="1101010111000100";
        when 5863 => y_in <= "10010110"; x_in <= "01100111"; z_correct<="1101010101011010";
        when 5864 => y_in <= "10010110"; x_in <= "01101000"; z_correct<="1101010011110000";
        when 5865 => y_in <= "10010110"; x_in <= "01101001"; z_correct<="1101010010000110";
        when 5866 => y_in <= "10010110"; x_in <= "01101010"; z_correct<="1101010000011100";
        when 5867 => y_in <= "10010110"; x_in <= "01101011"; z_correct<="1101001110110010";
        when 5868 => y_in <= "10010110"; x_in <= "01101100"; z_correct<="1101001101001000";
        when 5869 => y_in <= "10010110"; x_in <= "01101101"; z_correct<="1101001011011110";
        when 5870 => y_in <= "10010110"; x_in <= "01101110"; z_correct<="1101001001110100";
        when 5871 => y_in <= "10010110"; x_in <= "01101111"; z_correct<="1101001000001010";
        when 5872 => y_in <= "10010110"; x_in <= "01110000"; z_correct<="1101000110100000";
        when 5873 => y_in <= "10010110"; x_in <= "01110001"; z_correct<="1101000100110110";
        when 5874 => y_in <= "10010110"; x_in <= "01110010"; z_correct<="1101000011001100";
        when 5875 => y_in <= "10010110"; x_in <= "01110011"; z_correct<="1101000001100010";
        when 5876 => y_in <= "10010110"; x_in <= "01110100"; z_correct<="1100111111111000";
        when 5877 => y_in <= "10010110"; x_in <= "01110101"; z_correct<="1100111110001110";
        when 5878 => y_in <= "10010110"; x_in <= "01110110"; z_correct<="1100111100100100";
        when 5879 => y_in <= "10010110"; x_in <= "01110111"; z_correct<="1100111010111010";
        when 5880 => y_in <= "10010110"; x_in <= "01111000"; z_correct<="1100111001010000";
        when 5881 => y_in <= "10010110"; x_in <= "01111001"; z_correct<="1100110111100110";
        when 5882 => y_in <= "10010110"; x_in <= "01111010"; z_correct<="1100110101111100";
        when 5883 => y_in <= "10010110"; x_in <= "01111011"; z_correct<="1100110100010010";
        when 5884 => y_in <= "10010110"; x_in <= "01111100"; z_correct<="1100110010101000";
        when 5885 => y_in <= "10010110"; x_in <= "01111101"; z_correct<="1100110000111110";
        when 5886 => y_in <= "10010110"; x_in <= "01111110"; z_correct<="1100101111010100";
        when 5887 => y_in <= "10010110"; x_in <= "01111111"; z_correct<="1100101101101010";
        when 5888 => y_in <= "10010111"; x_in <= "10000000"; z_correct<="0011010010000000";
        when 5889 => y_in <= "10010111"; x_in <= "10000001"; z_correct<="0011010000010111";
        when 5890 => y_in <= "10010111"; x_in <= "10000010"; z_correct<="0011001110101110";
        when 5891 => y_in <= "10010111"; x_in <= "10000011"; z_correct<="0011001101000101";
        when 5892 => y_in <= "10010111"; x_in <= "10000100"; z_correct<="0011001011011100";
        when 5893 => y_in <= "10010111"; x_in <= "10000101"; z_correct<="0011001001110011";
        when 5894 => y_in <= "10010111"; x_in <= "10000110"; z_correct<="0011001000001010";
        when 5895 => y_in <= "10010111"; x_in <= "10000111"; z_correct<="0011000110100001";
        when 5896 => y_in <= "10010111"; x_in <= "10001000"; z_correct<="0011000100111000";
        when 5897 => y_in <= "10010111"; x_in <= "10001001"; z_correct<="0011000011001111";
        when 5898 => y_in <= "10010111"; x_in <= "10001010"; z_correct<="0011000001100110";
        when 5899 => y_in <= "10010111"; x_in <= "10001011"; z_correct<="0010111111111101";
        when 5900 => y_in <= "10010111"; x_in <= "10001100"; z_correct<="0010111110010100";
        when 5901 => y_in <= "10010111"; x_in <= "10001101"; z_correct<="0010111100101011";
        when 5902 => y_in <= "10010111"; x_in <= "10001110"; z_correct<="0010111011000010";
        when 5903 => y_in <= "10010111"; x_in <= "10001111"; z_correct<="0010111001011001";
        when 5904 => y_in <= "10010111"; x_in <= "10010000"; z_correct<="0010110111110000";
        when 5905 => y_in <= "10010111"; x_in <= "10010001"; z_correct<="0010110110000111";
        when 5906 => y_in <= "10010111"; x_in <= "10010010"; z_correct<="0010110100011110";
        when 5907 => y_in <= "10010111"; x_in <= "10010011"; z_correct<="0010110010110101";
        when 5908 => y_in <= "10010111"; x_in <= "10010100"; z_correct<="0010110001001100";
        when 5909 => y_in <= "10010111"; x_in <= "10010101"; z_correct<="0010101111100011";
        when 5910 => y_in <= "10010111"; x_in <= "10010110"; z_correct<="0010101101111010";
        when 5911 => y_in <= "10010111"; x_in <= "10010111"; z_correct<="0010101100010001";
        when 5912 => y_in <= "10010111"; x_in <= "10011000"; z_correct<="0010101010101000";
        when 5913 => y_in <= "10010111"; x_in <= "10011001"; z_correct<="0010101000111111";
        when 5914 => y_in <= "10010111"; x_in <= "10011010"; z_correct<="0010100111010110";
        when 5915 => y_in <= "10010111"; x_in <= "10011011"; z_correct<="0010100101101101";
        when 5916 => y_in <= "10010111"; x_in <= "10011100"; z_correct<="0010100100000100";
        when 5917 => y_in <= "10010111"; x_in <= "10011101"; z_correct<="0010100010011011";
        when 5918 => y_in <= "10010111"; x_in <= "10011110"; z_correct<="0010100000110010";
        when 5919 => y_in <= "10010111"; x_in <= "10011111"; z_correct<="0010011111001001";
        when 5920 => y_in <= "10010111"; x_in <= "10100000"; z_correct<="0010011101100000";
        when 5921 => y_in <= "10010111"; x_in <= "10100001"; z_correct<="0010011011110111";
        when 5922 => y_in <= "10010111"; x_in <= "10100010"; z_correct<="0010011010001110";
        when 5923 => y_in <= "10010111"; x_in <= "10100011"; z_correct<="0010011000100101";
        when 5924 => y_in <= "10010111"; x_in <= "10100100"; z_correct<="0010010110111100";
        when 5925 => y_in <= "10010111"; x_in <= "10100101"; z_correct<="0010010101010011";
        when 5926 => y_in <= "10010111"; x_in <= "10100110"; z_correct<="0010010011101010";
        when 5927 => y_in <= "10010111"; x_in <= "10100111"; z_correct<="0010010010000001";
        when 5928 => y_in <= "10010111"; x_in <= "10101000"; z_correct<="0010010000011000";
        when 5929 => y_in <= "10010111"; x_in <= "10101001"; z_correct<="0010001110101111";
        when 5930 => y_in <= "10010111"; x_in <= "10101010"; z_correct<="0010001101000110";
        when 5931 => y_in <= "10010111"; x_in <= "10101011"; z_correct<="0010001011011101";
        when 5932 => y_in <= "10010111"; x_in <= "10101100"; z_correct<="0010001001110100";
        when 5933 => y_in <= "10010111"; x_in <= "10101101"; z_correct<="0010001000001011";
        when 5934 => y_in <= "10010111"; x_in <= "10101110"; z_correct<="0010000110100010";
        when 5935 => y_in <= "10010111"; x_in <= "10101111"; z_correct<="0010000100111001";
        when 5936 => y_in <= "10010111"; x_in <= "10110000"; z_correct<="0010000011010000";
        when 5937 => y_in <= "10010111"; x_in <= "10110001"; z_correct<="0010000001100111";
        when 5938 => y_in <= "10010111"; x_in <= "10110010"; z_correct<="0001111111111110";
        when 5939 => y_in <= "10010111"; x_in <= "10110011"; z_correct<="0001111110010101";
        when 5940 => y_in <= "10010111"; x_in <= "10110100"; z_correct<="0001111100101100";
        when 5941 => y_in <= "10010111"; x_in <= "10110101"; z_correct<="0001111011000011";
        when 5942 => y_in <= "10010111"; x_in <= "10110110"; z_correct<="0001111001011010";
        when 5943 => y_in <= "10010111"; x_in <= "10110111"; z_correct<="0001110111110001";
        when 5944 => y_in <= "10010111"; x_in <= "10111000"; z_correct<="0001110110001000";
        when 5945 => y_in <= "10010111"; x_in <= "10111001"; z_correct<="0001110100011111";
        when 5946 => y_in <= "10010111"; x_in <= "10111010"; z_correct<="0001110010110110";
        when 5947 => y_in <= "10010111"; x_in <= "10111011"; z_correct<="0001110001001101";
        when 5948 => y_in <= "10010111"; x_in <= "10111100"; z_correct<="0001101111100100";
        when 5949 => y_in <= "10010111"; x_in <= "10111101"; z_correct<="0001101101111011";
        when 5950 => y_in <= "10010111"; x_in <= "10111110"; z_correct<="0001101100010010";
        when 5951 => y_in <= "10010111"; x_in <= "10111111"; z_correct<="0001101010101001";
        when 5952 => y_in <= "10010111"; x_in <= "11000000"; z_correct<="0001101001000000";
        when 5953 => y_in <= "10010111"; x_in <= "11000001"; z_correct<="0001100111010111";
        when 5954 => y_in <= "10010111"; x_in <= "11000010"; z_correct<="0001100101101110";
        when 5955 => y_in <= "10010111"; x_in <= "11000011"; z_correct<="0001100100000101";
        when 5956 => y_in <= "10010111"; x_in <= "11000100"; z_correct<="0001100010011100";
        when 5957 => y_in <= "10010111"; x_in <= "11000101"; z_correct<="0001100000110011";
        when 5958 => y_in <= "10010111"; x_in <= "11000110"; z_correct<="0001011111001010";
        when 5959 => y_in <= "10010111"; x_in <= "11000111"; z_correct<="0001011101100001";
        when 5960 => y_in <= "10010111"; x_in <= "11001000"; z_correct<="0001011011111000";
        when 5961 => y_in <= "10010111"; x_in <= "11001001"; z_correct<="0001011010001111";
        when 5962 => y_in <= "10010111"; x_in <= "11001010"; z_correct<="0001011000100110";
        when 5963 => y_in <= "10010111"; x_in <= "11001011"; z_correct<="0001010110111101";
        when 5964 => y_in <= "10010111"; x_in <= "11001100"; z_correct<="0001010101010100";
        when 5965 => y_in <= "10010111"; x_in <= "11001101"; z_correct<="0001010011101011";
        when 5966 => y_in <= "10010111"; x_in <= "11001110"; z_correct<="0001010010000010";
        when 5967 => y_in <= "10010111"; x_in <= "11001111"; z_correct<="0001010000011001";
        when 5968 => y_in <= "10010111"; x_in <= "11010000"; z_correct<="0001001110110000";
        when 5969 => y_in <= "10010111"; x_in <= "11010001"; z_correct<="0001001101000111";
        when 5970 => y_in <= "10010111"; x_in <= "11010010"; z_correct<="0001001011011110";
        when 5971 => y_in <= "10010111"; x_in <= "11010011"; z_correct<="0001001001110101";
        when 5972 => y_in <= "10010111"; x_in <= "11010100"; z_correct<="0001001000001100";
        when 5973 => y_in <= "10010111"; x_in <= "11010101"; z_correct<="0001000110100011";
        when 5974 => y_in <= "10010111"; x_in <= "11010110"; z_correct<="0001000100111010";
        when 5975 => y_in <= "10010111"; x_in <= "11010111"; z_correct<="0001000011010001";
        when 5976 => y_in <= "10010111"; x_in <= "11011000"; z_correct<="0001000001101000";
        when 5977 => y_in <= "10010111"; x_in <= "11011001"; z_correct<="0000111111111111";
        when 5978 => y_in <= "10010111"; x_in <= "11011010"; z_correct<="0000111110010110";
        when 5979 => y_in <= "10010111"; x_in <= "11011011"; z_correct<="0000111100101101";
        when 5980 => y_in <= "10010111"; x_in <= "11011100"; z_correct<="0000111011000100";
        when 5981 => y_in <= "10010111"; x_in <= "11011101"; z_correct<="0000111001011011";
        when 5982 => y_in <= "10010111"; x_in <= "11011110"; z_correct<="0000110111110010";
        when 5983 => y_in <= "10010111"; x_in <= "11011111"; z_correct<="0000110110001001";
        when 5984 => y_in <= "10010111"; x_in <= "11100000"; z_correct<="0000110100100000";
        when 5985 => y_in <= "10010111"; x_in <= "11100001"; z_correct<="0000110010110111";
        when 5986 => y_in <= "10010111"; x_in <= "11100010"; z_correct<="0000110001001110";
        when 5987 => y_in <= "10010111"; x_in <= "11100011"; z_correct<="0000101111100101";
        when 5988 => y_in <= "10010111"; x_in <= "11100100"; z_correct<="0000101101111100";
        when 5989 => y_in <= "10010111"; x_in <= "11100101"; z_correct<="0000101100010011";
        when 5990 => y_in <= "10010111"; x_in <= "11100110"; z_correct<="0000101010101010";
        when 5991 => y_in <= "10010111"; x_in <= "11100111"; z_correct<="0000101001000001";
        when 5992 => y_in <= "10010111"; x_in <= "11101000"; z_correct<="0000100111011000";
        when 5993 => y_in <= "10010111"; x_in <= "11101001"; z_correct<="0000100101101111";
        when 5994 => y_in <= "10010111"; x_in <= "11101010"; z_correct<="0000100100000110";
        when 5995 => y_in <= "10010111"; x_in <= "11101011"; z_correct<="0000100010011101";
        when 5996 => y_in <= "10010111"; x_in <= "11101100"; z_correct<="0000100000110100";
        when 5997 => y_in <= "10010111"; x_in <= "11101101"; z_correct<="0000011111001011";
        when 5998 => y_in <= "10010111"; x_in <= "11101110"; z_correct<="0000011101100010";
        when 5999 => y_in <= "10010111"; x_in <= "11101111"; z_correct<="0000011011111001";
        when 6000 => y_in <= "10010111"; x_in <= "11110000"; z_correct<="0000011010010000";
        when 6001 => y_in <= "10010111"; x_in <= "11110001"; z_correct<="0000011000100111";
        when 6002 => y_in <= "10010111"; x_in <= "11110010"; z_correct<="0000010110111110";
        when 6003 => y_in <= "10010111"; x_in <= "11110011"; z_correct<="0000010101010101";
        when 6004 => y_in <= "10010111"; x_in <= "11110100"; z_correct<="0000010011101100";
        when 6005 => y_in <= "10010111"; x_in <= "11110101"; z_correct<="0000010010000011";
        when 6006 => y_in <= "10010111"; x_in <= "11110110"; z_correct<="0000010000011010";
        when 6007 => y_in <= "10010111"; x_in <= "11110111"; z_correct<="0000001110110001";
        when 6008 => y_in <= "10010111"; x_in <= "11111000"; z_correct<="0000001101001000";
        when 6009 => y_in <= "10010111"; x_in <= "11111001"; z_correct<="0000001011011111";
        when 6010 => y_in <= "10010111"; x_in <= "11111010"; z_correct<="0000001001110110";
        when 6011 => y_in <= "10010111"; x_in <= "11111011"; z_correct<="0000001000001101";
        when 6012 => y_in <= "10010111"; x_in <= "11111100"; z_correct<="0000000110100100";
        when 6013 => y_in <= "10010111"; x_in <= "11111101"; z_correct<="0000000100111011";
        when 6014 => y_in <= "10010111"; x_in <= "11111110"; z_correct<="0000000011010010";
        when 6015 => y_in <= "10010111"; x_in <= "11111111"; z_correct<="0000000001101001";
        when 6016 => y_in <= "10010111"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 6017 => y_in <= "10010111"; x_in <= "00000001"; z_correct<="1111111110010111";
        when 6018 => y_in <= "10010111"; x_in <= "00000010"; z_correct<="1111111100101110";
        when 6019 => y_in <= "10010111"; x_in <= "00000011"; z_correct<="1111111011000101";
        when 6020 => y_in <= "10010111"; x_in <= "00000100"; z_correct<="1111111001011100";
        when 6021 => y_in <= "10010111"; x_in <= "00000101"; z_correct<="1111110111110011";
        when 6022 => y_in <= "10010111"; x_in <= "00000110"; z_correct<="1111110110001010";
        when 6023 => y_in <= "10010111"; x_in <= "00000111"; z_correct<="1111110100100001";
        when 6024 => y_in <= "10010111"; x_in <= "00001000"; z_correct<="1111110010111000";
        when 6025 => y_in <= "10010111"; x_in <= "00001001"; z_correct<="1111110001001111";
        when 6026 => y_in <= "10010111"; x_in <= "00001010"; z_correct<="1111101111100110";
        when 6027 => y_in <= "10010111"; x_in <= "00001011"; z_correct<="1111101101111101";
        when 6028 => y_in <= "10010111"; x_in <= "00001100"; z_correct<="1111101100010100";
        when 6029 => y_in <= "10010111"; x_in <= "00001101"; z_correct<="1111101010101011";
        when 6030 => y_in <= "10010111"; x_in <= "00001110"; z_correct<="1111101001000010";
        when 6031 => y_in <= "10010111"; x_in <= "00001111"; z_correct<="1111100111011001";
        when 6032 => y_in <= "10010111"; x_in <= "00010000"; z_correct<="1111100101110000";
        when 6033 => y_in <= "10010111"; x_in <= "00010001"; z_correct<="1111100100000111";
        when 6034 => y_in <= "10010111"; x_in <= "00010010"; z_correct<="1111100010011110";
        when 6035 => y_in <= "10010111"; x_in <= "00010011"; z_correct<="1111100000110101";
        when 6036 => y_in <= "10010111"; x_in <= "00010100"; z_correct<="1111011111001100";
        when 6037 => y_in <= "10010111"; x_in <= "00010101"; z_correct<="1111011101100011";
        when 6038 => y_in <= "10010111"; x_in <= "00010110"; z_correct<="1111011011111010";
        when 6039 => y_in <= "10010111"; x_in <= "00010111"; z_correct<="1111011010010001";
        when 6040 => y_in <= "10010111"; x_in <= "00011000"; z_correct<="1111011000101000";
        when 6041 => y_in <= "10010111"; x_in <= "00011001"; z_correct<="1111010110111111";
        when 6042 => y_in <= "10010111"; x_in <= "00011010"; z_correct<="1111010101010110";
        when 6043 => y_in <= "10010111"; x_in <= "00011011"; z_correct<="1111010011101101";
        when 6044 => y_in <= "10010111"; x_in <= "00011100"; z_correct<="1111010010000100";
        when 6045 => y_in <= "10010111"; x_in <= "00011101"; z_correct<="1111010000011011";
        when 6046 => y_in <= "10010111"; x_in <= "00011110"; z_correct<="1111001110110010";
        when 6047 => y_in <= "10010111"; x_in <= "00011111"; z_correct<="1111001101001001";
        when 6048 => y_in <= "10010111"; x_in <= "00100000"; z_correct<="1111001011100000";
        when 6049 => y_in <= "10010111"; x_in <= "00100001"; z_correct<="1111001001110111";
        when 6050 => y_in <= "10010111"; x_in <= "00100010"; z_correct<="1111001000001110";
        when 6051 => y_in <= "10010111"; x_in <= "00100011"; z_correct<="1111000110100101";
        when 6052 => y_in <= "10010111"; x_in <= "00100100"; z_correct<="1111000100111100";
        when 6053 => y_in <= "10010111"; x_in <= "00100101"; z_correct<="1111000011010011";
        when 6054 => y_in <= "10010111"; x_in <= "00100110"; z_correct<="1111000001101010";
        when 6055 => y_in <= "10010111"; x_in <= "00100111"; z_correct<="1111000000000001";
        when 6056 => y_in <= "10010111"; x_in <= "00101000"; z_correct<="1110111110011000";
        when 6057 => y_in <= "10010111"; x_in <= "00101001"; z_correct<="1110111100101111";
        when 6058 => y_in <= "10010111"; x_in <= "00101010"; z_correct<="1110111011000110";
        when 6059 => y_in <= "10010111"; x_in <= "00101011"; z_correct<="1110111001011101";
        when 6060 => y_in <= "10010111"; x_in <= "00101100"; z_correct<="1110110111110100";
        when 6061 => y_in <= "10010111"; x_in <= "00101101"; z_correct<="1110110110001011";
        when 6062 => y_in <= "10010111"; x_in <= "00101110"; z_correct<="1110110100100010";
        when 6063 => y_in <= "10010111"; x_in <= "00101111"; z_correct<="1110110010111001";
        when 6064 => y_in <= "10010111"; x_in <= "00110000"; z_correct<="1110110001010000";
        when 6065 => y_in <= "10010111"; x_in <= "00110001"; z_correct<="1110101111100111";
        when 6066 => y_in <= "10010111"; x_in <= "00110010"; z_correct<="1110101101111110";
        when 6067 => y_in <= "10010111"; x_in <= "00110011"; z_correct<="1110101100010101";
        when 6068 => y_in <= "10010111"; x_in <= "00110100"; z_correct<="1110101010101100";
        when 6069 => y_in <= "10010111"; x_in <= "00110101"; z_correct<="1110101001000011";
        when 6070 => y_in <= "10010111"; x_in <= "00110110"; z_correct<="1110100111011010";
        when 6071 => y_in <= "10010111"; x_in <= "00110111"; z_correct<="1110100101110001";
        when 6072 => y_in <= "10010111"; x_in <= "00111000"; z_correct<="1110100100001000";
        when 6073 => y_in <= "10010111"; x_in <= "00111001"; z_correct<="1110100010011111";
        when 6074 => y_in <= "10010111"; x_in <= "00111010"; z_correct<="1110100000110110";
        when 6075 => y_in <= "10010111"; x_in <= "00111011"; z_correct<="1110011111001101";
        when 6076 => y_in <= "10010111"; x_in <= "00111100"; z_correct<="1110011101100100";
        when 6077 => y_in <= "10010111"; x_in <= "00111101"; z_correct<="1110011011111011";
        when 6078 => y_in <= "10010111"; x_in <= "00111110"; z_correct<="1110011010010010";
        when 6079 => y_in <= "10010111"; x_in <= "00111111"; z_correct<="1110011000101001";
        when 6080 => y_in <= "10010111"; x_in <= "01000000"; z_correct<="1110010111000000";
        when 6081 => y_in <= "10010111"; x_in <= "01000001"; z_correct<="1110010101010111";
        when 6082 => y_in <= "10010111"; x_in <= "01000010"; z_correct<="1110010011101110";
        when 6083 => y_in <= "10010111"; x_in <= "01000011"; z_correct<="1110010010000101";
        when 6084 => y_in <= "10010111"; x_in <= "01000100"; z_correct<="1110010000011100";
        when 6085 => y_in <= "10010111"; x_in <= "01000101"; z_correct<="1110001110110011";
        when 6086 => y_in <= "10010111"; x_in <= "01000110"; z_correct<="1110001101001010";
        when 6087 => y_in <= "10010111"; x_in <= "01000111"; z_correct<="1110001011100001";
        when 6088 => y_in <= "10010111"; x_in <= "01001000"; z_correct<="1110001001111000";
        when 6089 => y_in <= "10010111"; x_in <= "01001001"; z_correct<="1110001000001111";
        when 6090 => y_in <= "10010111"; x_in <= "01001010"; z_correct<="1110000110100110";
        when 6091 => y_in <= "10010111"; x_in <= "01001011"; z_correct<="1110000100111101";
        when 6092 => y_in <= "10010111"; x_in <= "01001100"; z_correct<="1110000011010100";
        when 6093 => y_in <= "10010111"; x_in <= "01001101"; z_correct<="1110000001101011";
        when 6094 => y_in <= "10010111"; x_in <= "01001110"; z_correct<="1110000000000010";
        when 6095 => y_in <= "10010111"; x_in <= "01001111"; z_correct<="1101111110011001";
        when 6096 => y_in <= "10010111"; x_in <= "01010000"; z_correct<="1101111100110000";
        when 6097 => y_in <= "10010111"; x_in <= "01010001"; z_correct<="1101111011000111";
        when 6098 => y_in <= "10010111"; x_in <= "01010010"; z_correct<="1101111001011110";
        when 6099 => y_in <= "10010111"; x_in <= "01010011"; z_correct<="1101110111110101";
        when 6100 => y_in <= "10010111"; x_in <= "01010100"; z_correct<="1101110110001100";
        when 6101 => y_in <= "10010111"; x_in <= "01010101"; z_correct<="1101110100100011";
        when 6102 => y_in <= "10010111"; x_in <= "01010110"; z_correct<="1101110010111010";
        when 6103 => y_in <= "10010111"; x_in <= "01010111"; z_correct<="1101110001010001";
        when 6104 => y_in <= "10010111"; x_in <= "01011000"; z_correct<="1101101111101000";
        when 6105 => y_in <= "10010111"; x_in <= "01011001"; z_correct<="1101101101111111";
        when 6106 => y_in <= "10010111"; x_in <= "01011010"; z_correct<="1101101100010110";
        when 6107 => y_in <= "10010111"; x_in <= "01011011"; z_correct<="1101101010101101";
        when 6108 => y_in <= "10010111"; x_in <= "01011100"; z_correct<="1101101001000100";
        when 6109 => y_in <= "10010111"; x_in <= "01011101"; z_correct<="1101100111011011";
        when 6110 => y_in <= "10010111"; x_in <= "01011110"; z_correct<="1101100101110010";
        when 6111 => y_in <= "10010111"; x_in <= "01011111"; z_correct<="1101100100001001";
        when 6112 => y_in <= "10010111"; x_in <= "01100000"; z_correct<="1101100010100000";
        when 6113 => y_in <= "10010111"; x_in <= "01100001"; z_correct<="1101100000110111";
        when 6114 => y_in <= "10010111"; x_in <= "01100010"; z_correct<="1101011111001110";
        when 6115 => y_in <= "10010111"; x_in <= "01100011"; z_correct<="1101011101100101";
        when 6116 => y_in <= "10010111"; x_in <= "01100100"; z_correct<="1101011011111100";
        when 6117 => y_in <= "10010111"; x_in <= "01100101"; z_correct<="1101011010010011";
        when 6118 => y_in <= "10010111"; x_in <= "01100110"; z_correct<="1101011000101010";
        when 6119 => y_in <= "10010111"; x_in <= "01100111"; z_correct<="1101010111000001";
        when 6120 => y_in <= "10010111"; x_in <= "01101000"; z_correct<="1101010101011000";
        when 6121 => y_in <= "10010111"; x_in <= "01101001"; z_correct<="1101010011101111";
        when 6122 => y_in <= "10010111"; x_in <= "01101010"; z_correct<="1101010010000110";
        when 6123 => y_in <= "10010111"; x_in <= "01101011"; z_correct<="1101010000011101";
        when 6124 => y_in <= "10010111"; x_in <= "01101100"; z_correct<="1101001110110100";
        when 6125 => y_in <= "10010111"; x_in <= "01101101"; z_correct<="1101001101001011";
        when 6126 => y_in <= "10010111"; x_in <= "01101110"; z_correct<="1101001011100010";
        when 6127 => y_in <= "10010111"; x_in <= "01101111"; z_correct<="1101001001111001";
        when 6128 => y_in <= "10010111"; x_in <= "01110000"; z_correct<="1101001000010000";
        when 6129 => y_in <= "10010111"; x_in <= "01110001"; z_correct<="1101000110100111";
        when 6130 => y_in <= "10010111"; x_in <= "01110010"; z_correct<="1101000100111110";
        when 6131 => y_in <= "10010111"; x_in <= "01110011"; z_correct<="1101000011010101";
        when 6132 => y_in <= "10010111"; x_in <= "01110100"; z_correct<="1101000001101100";
        when 6133 => y_in <= "10010111"; x_in <= "01110101"; z_correct<="1101000000000011";
        when 6134 => y_in <= "10010111"; x_in <= "01110110"; z_correct<="1100111110011010";
        when 6135 => y_in <= "10010111"; x_in <= "01110111"; z_correct<="1100111100110001";
        when 6136 => y_in <= "10010111"; x_in <= "01111000"; z_correct<="1100111011001000";
        when 6137 => y_in <= "10010111"; x_in <= "01111001"; z_correct<="1100111001011111";
        when 6138 => y_in <= "10010111"; x_in <= "01111010"; z_correct<="1100110111110110";
        when 6139 => y_in <= "10010111"; x_in <= "01111011"; z_correct<="1100110110001101";
        when 6140 => y_in <= "10010111"; x_in <= "01111100"; z_correct<="1100110100100100";
        when 6141 => y_in <= "10010111"; x_in <= "01111101"; z_correct<="1100110010111011";
        when 6142 => y_in <= "10010111"; x_in <= "01111110"; z_correct<="1100110001010010";
        when 6143 => y_in <= "10010111"; x_in <= "01111111"; z_correct<="1100101111101001";
        when 6144 => y_in <= "10011000"; x_in <= "10000000"; z_correct<="0011010000000000";
        when 6145 => y_in <= "10011000"; x_in <= "10000001"; z_correct<="0011001110011000";
        when 6146 => y_in <= "10011000"; x_in <= "10000010"; z_correct<="0011001100110000";
        when 6147 => y_in <= "10011000"; x_in <= "10000011"; z_correct<="0011001011001000";
        when 6148 => y_in <= "10011000"; x_in <= "10000100"; z_correct<="0011001001100000";
        when 6149 => y_in <= "10011000"; x_in <= "10000101"; z_correct<="0011000111111000";
        when 6150 => y_in <= "10011000"; x_in <= "10000110"; z_correct<="0011000110010000";
        when 6151 => y_in <= "10011000"; x_in <= "10000111"; z_correct<="0011000100101000";
        when 6152 => y_in <= "10011000"; x_in <= "10001000"; z_correct<="0011000011000000";
        when 6153 => y_in <= "10011000"; x_in <= "10001001"; z_correct<="0011000001011000";
        when 6154 => y_in <= "10011000"; x_in <= "10001010"; z_correct<="0010111111110000";
        when 6155 => y_in <= "10011000"; x_in <= "10001011"; z_correct<="0010111110001000";
        when 6156 => y_in <= "10011000"; x_in <= "10001100"; z_correct<="0010111100100000";
        when 6157 => y_in <= "10011000"; x_in <= "10001101"; z_correct<="0010111010111000";
        when 6158 => y_in <= "10011000"; x_in <= "10001110"; z_correct<="0010111001010000";
        when 6159 => y_in <= "10011000"; x_in <= "10001111"; z_correct<="0010110111101000";
        when 6160 => y_in <= "10011000"; x_in <= "10010000"; z_correct<="0010110110000000";
        when 6161 => y_in <= "10011000"; x_in <= "10010001"; z_correct<="0010110100011000";
        when 6162 => y_in <= "10011000"; x_in <= "10010010"; z_correct<="0010110010110000";
        when 6163 => y_in <= "10011000"; x_in <= "10010011"; z_correct<="0010110001001000";
        when 6164 => y_in <= "10011000"; x_in <= "10010100"; z_correct<="0010101111100000";
        when 6165 => y_in <= "10011000"; x_in <= "10010101"; z_correct<="0010101101111000";
        when 6166 => y_in <= "10011000"; x_in <= "10010110"; z_correct<="0010101100010000";
        when 6167 => y_in <= "10011000"; x_in <= "10010111"; z_correct<="0010101010101000";
        when 6168 => y_in <= "10011000"; x_in <= "10011000"; z_correct<="0010101001000000";
        when 6169 => y_in <= "10011000"; x_in <= "10011001"; z_correct<="0010100111011000";
        when 6170 => y_in <= "10011000"; x_in <= "10011010"; z_correct<="0010100101110000";
        when 6171 => y_in <= "10011000"; x_in <= "10011011"; z_correct<="0010100100001000";
        when 6172 => y_in <= "10011000"; x_in <= "10011100"; z_correct<="0010100010100000";
        when 6173 => y_in <= "10011000"; x_in <= "10011101"; z_correct<="0010100000111000";
        when 6174 => y_in <= "10011000"; x_in <= "10011110"; z_correct<="0010011111010000";
        when 6175 => y_in <= "10011000"; x_in <= "10011111"; z_correct<="0010011101101000";
        when 6176 => y_in <= "10011000"; x_in <= "10100000"; z_correct<="0010011100000000";
        when 6177 => y_in <= "10011000"; x_in <= "10100001"; z_correct<="0010011010011000";
        when 6178 => y_in <= "10011000"; x_in <= "10100010"; z_correct<="0010011000110000";
        when 6179 => y_in <= "10011000"; x_in <= "10100011"; z_correct<="0010010111001000";
        when 6180 => y_in <= "10011000"; x_in <= "10100100"; z_correct<="0010010101100000";
        when 6181 => y_in <= "10011000"; x_in <= "10100101"; z_correct<="0010010011111000";
        when 6182 => y_in <= "10011000"; x_in <= "10100110"; z_correct<="0010010010010000";
        when 6183 => y_in <= "10011000"; x_in <= "10100111"; z_correct<="0010010000101000";
        when 6184 => y_in <= "10011000"; x_in <= "10101000"; z_correct<="0010001111000000";
        when 6185 => y_in <= "10011000"; x_in <= "10101001"; z_correct<="0010001101011000";
        when 6186 => y_in <= "10011000"; x_in <= "10101010"; z_correct<="0010001011110000";
        when 6187 => y_in <= "10011000"; x_in <= "10101011"; z_correct<="0010001010001000";
        when 6188 => y_in <= "10011000"; x_in <= "10101100"; z_correct<="0010001000100000";
        when 6189 => y_in <= "10011000"; x_in <= "10101101"; z_correct<="0010000110111000";
        when 6190 => y_in <= "10011000"; x_in <= "10101110"; z_correct<="0010000101010000";
        when 6191 => y_in <= "10011000"; x_in <= "10101111"; z_correct<="0010000011101000";
        when 6192 => y_in <= "10011000"; x_in <= "10110000"; z_correct<="0010000010000000";
        when 6193 => y_in <= "10011000"; x_in <= "10110001"; z_correct<="0010000000011000";
        when 6194 => y_in <= "10011000"; x_in <= "10110010"; z_correct<="0001111110110000";
        when 6195 => y_in <= "10011000"; x_in <= "10110011"; z_correct<="0001111101001000";
        when 6196 => y_in <= "10011000"; x_in <= "10110100"; z_correct<="0001111011100000";
        when 6197 => y_in <= "10011000"; x_in <= "10110101"; z_correct<="0001111001111000";
        when 6198 => y_in <= "10011000"; x_in <= "10110110"; z_correct<="0001111000010000";
        when 6199 => y_in <= "10011000"; x_in <= "10110111"; z_correct<="0001110110101000";
        when 6200 => y_in <= "10011000"; x_in <= "10111000"; z_correct<="0001110101000000";
        when 6201 => y_in <= "10011000"; x_in <= "10111001"; z_correct<="0001110011011000";
        when 6202 => y_in <= "10011000"; x_in <= "10111010"; z_correct<="0001110001110000";
        when 6203 => y_in <= "10011000"; x_in <= "10111011"; z_correct<="0001110000001000";
        when 6204 => y_in <= "10011000"; x_in <= "10111100"; z_correct<="0001101110100000";
        when 6205 => y_in <= "10011000"; x_in <= "10111101"; z_correct<="0001101100111000";
        when 6206 => y_in <= "10011000"; x_in <= "10111110"; z_correct<="0001101011010000";
        when 6207 => y_in <= "10011000"; x_in <= "10111111"; z_correct<="0001101001101000";
        when 6208 => y_in <= "10011000"; x_in <= "11000000"; z_correct<="0001101000000000";
        when 6209 => y_in <= "10011000"; x_in <= "11000001"; z_correct<="0001100110011000";
        when 6210 => y_in <= "10011000"; x_in <= "11000010"; z_correct<="0001100100110000";
        when 6211 => y_in <= "10011000"; x_in <= "11000011"; z_correct<="0001100011001000";
        when 6212 => y_in <= "10011000"; x_in <= "11000100"; z_correct<="0001100001100000";
        when 6213 => y_in <= "10011000"; x_in <= "11000101"; z_correct<="0001011111111000";
        when 6214 => y_in <= "10011000"; x_in <= "11000110"; z_correct<="0001011110010000";
        when 6215 => y_in <= "10011000"; x_in <= "11000111"; z_correct<="0001011100101000";
        when 6216 => y_in <= "10011000"; x_in <= "11001000"; z_correct<="0001011011000000";
        when 6217 => y_in <= "10011000"; x_in <= "11001001"; z_correct<="0001011001011000";
        when 6218 => y_in <= "10011000"; x_in <= "11001010"; z_correct<="0001010111110000";
        when 6219 => y_in <= "10011000"; x_in <= "11001011"; z_correct<="0001010110001000";
        when 6220 => y_in <= "10011000"; x_in <= "11001100"; z_correct<="0001010100100000";
        when 6221 => y_in <= "10011000"; x_in <= "11001101"; z_correct<="0001010010111000";
        when 6222 => y_in <= "10011000"; x_in <= "11001110"; z_correct<="0001010001010000";
        when 6223 => y_in <= "10011000"; x_in <= "11001111"; z_correct<="0001001111101000";
        when 6224 => y_in <= "10011000"; x_in <= "11010000"; z_correct<="0001001110000000";
        when 6225 => y_in <= "10011000"; x_in <= "11010001"; z_correct<="0001001100011000";
        when 6226 => y_in <= "10011000"; x_in <= "11010010"; z_correct<="0001001010110000";
        when 6227 => y_in <= "10011000"; x_in <= "11010011"; z_correct<="0001001001001000";
        when 6228 => y_in <= "10011000"; x_in <= "11010100"; z_correct<="0001000111100000";
        when 6229 => y_in <= "10011000"; x_in <= "11010101"; z_correct<="0001000101111000";
        when 6230 => y_in <= "10011000"; x_in <= "11010110"; z_correct<="0001000100010000";
        when 6231 => y_in <= "10011000"; x_in <= "11010111"; z_correct<="0001000010101000";
        when 6232 => y_in <= "10011000"; x_in <= "11011000"; z_correct<="0001000001000000";
        when 6233 => y_in <= "10011000"; x_in <= "11011001"; z_correct<="0000111111011000";
        when 6234 => y_in <= "10011000"; x_in <= "11011010"; z_correct<="0000111101110000";
        when 6235 => y_in <= "10011000"; x_in <= "11011011"; z_correct<="0000111100001000";
        when 6236 => y_in <= "10011000"; x_in <= "11011100"; z_correct<="0000111010100000";
        when 6237 => y_in <= "10011000"; x_in <= "11011101"; z_correct<="0000111000111000";
        when 6238 => y_in <= "10011000"; x_in <= "11011110"; z_correct<="0000110111010000";
        when 6239 => y_in <= "10011000"; x_in <= "11011111"; z_correct<="0000110101101000";
        when 6240 => y_in <= "10011000"; x_in <= "11100000"; z_correct<="0000110100000000";
        when 6241 => y_in <= "10011000"; x_in <= "11100001"; z_correct<="0000110010011000";
        when 6242 => y_in <= "10011000"; x_in <= "11100010"; z_correct<="0000110000110000";
        when 6243 => y_in <= "10011000"; x_in <= "11100011"; z_correct<="0000101111001000";
        when 6244 => y_in <= "10011000"; x_in <= "11100100"; z_correct<="0000101101100000";
        when 6245 => y_in <= "10011000"; x_in <= "11100101"; z_correct<="0000101011111000";
        when 6246 => y_in <= "10011000"; x_in <= "11100110"; z_correct<="0000101010010000";
        when 6247 => y_in <= "10011000"; x_in <= "11100111"; z_correct<="0000101000101000";
        when 6248 => y_in <= "10011000"; x_in <= "11101000"; z_correct<="0000100111000000";
        when 6249 => y_in <= "10011000"; x_in <= "11101001"; z_correct<="0000100101011000";
        when 6250 => y_in <= "10011000"; x_in <= "11101010"; z_correct<="0000100011110000";
        when 6251 => y_in <= "10011000"; x_in <= "11101011"; z_correct<="0000100010001000";
        when 6252 => y_in <= "10011000"; x_in <= "11101100"; z_correct<="0000100000100000";
        when 6253 => y_in <= "10011000"; x_in <= "11101101"; z_correct<="0000011110111000";
        when 6254 => y_in <= "10011000"; x_in <= "11101110"; z_correct<="0000011101010000";
        when 6255 => y_in <= "10011000"; x_in <= "11101111"; z_correct<="0000011011101000";
        when 6256 => y_in <= "10011000"; x_in <= "11110000"; z_correct<="0000011010000000";
        when 6257 => y_in <= "10011000"; x_in <= "11110001"; z_correct<="0000011000011000";
        when 6258 => y_in <= "10011000"; x_in <= "11110010"; z_correct<="0000010110110000";
        when 6259 => y_in <= "10011000"; x_in <= "11110011"; z_correct<="0000010101001000";
        when 6260 => y_in <= "10011000"; x_in <= "11110100"; z_correct<="0000010011100000";
        when 6261 => y_in <= "10011000"; x_in <= "11110101"; z_correct<="0000010001111000";
        when 6262 => y_in <= "10011000"; x_in <= "11110110"; z_correct<="0000010000010000";
        when 6263 => y_in <= "10011000"; x_in <= "11110111"; z_correct<="0000001110101000";
        when 6264 => y_in <= "10011000"; x_in <= "11111000"; z_correct<="0000001101000000";
        when 6265 => y_in <= "10011000"; x_in <= "11111001"; z_correct<="0000001011011000";
        when 6266 => y_in <= "10011000"; x_in <= "11111010"; z_correct<="0000001001110000";
        when 6267 => y_in <= "10011000"; x_in <= "11111011"; z_correct<="0000001000001000";
        when 6268 => y_in <= "10011000"; x_in <= "11111100"; z_correct<="0000000110100000";
        when 6269 => y_in <= "10011000"; x_in <= "11111101"; z_correct<="0000000100111000";
        when 6270 => y_in <= "10011000"; x_in <= "11111110"; z_correct<="0000000011010000";
        when 6271 => y_in <= "10011000"; x_in <= "11111111"; z_correct<="0000000001101000";
        when 6272 => y_in <= "10011000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 6273 => y_in <= "10011000"; x_in <= "00000001"; z_correct<="1111111110011000";
        when 6274 => y_in <= "10011000"; x_in <= "00000010"; z_correct<="1111111100110000";
        when 6275 => y_in <= "10011000"; x_in <= "00000011"; z_correct<="1111111011001000";
        when 6276 => y_in <= "10011000"; x_in <= "00000100"; z_correct<="1111111001100000";
        when 6277 => y_in <= "10011000"; x_in <= "00000101"; z_correct<="1111110111111000";
        when 6278 => y_in <= "10011000"; x_in <= "00000110"; z_correct<="1111110110010000";
        when 6279 => y_in <= "10011000"; x_in <= "00000111"; z_correct<="1111110100101000";
        when 6280 => y_in <= "10011000"; x_in <= "00001000"; z_correct<="1111110011000000";
        when 6281 => y_in <= "10011000"; x_in <= "00001001"; z_correct<="1111110001011000";
        when 6282 => y_in <= "10011000"; x_in <= "00001010"; z_correct<="1111101111110000";
        when 6283 => y_in <= "10011000"; x_in <= "00001011"; z_correct<="1111101110001000";
        when 6284 => y_in <= "10011000"; x_in <= "00001100"; z_correct<="1111101100100000";
        when 6285 => y_in <= "10011000"; x_in <= "00001101"; z_correct<="1111101010111000";
        when 6286 => y_in <= "10011000"; x_in <= "00001110"; z_correct<="1111101001010000";
        when 6287 => y_in <= "10011000"; x_in <= "00001111"; z_correct<="1111100111101000";
        when 6288 => y_in <= "10011000"; x_in <= "00010000"; z_correct<="1111100110000000";
        when 6289 => y_in <= "10011000"; x_in <= "00010001"; z_correct<="1111100100011000";
        when 6290 => y_in <= "10011000"; x_in <= "00010010"; z_correct<="1111100010110000";
        when 6291 => y_in <= "10011000"; x_in <= "00010011"; z_correct<="1111100001001000";
        when 6292 => y_in <= "10011000"; x_in <= "00010100"; z_correct<="1111011111100000";
        when 6293 => y_in <= "10011000"; x_in <= "00010101"; z_correct<="1111011101111000";
        when 6294 => y_in <= "10011000"; x_in <= "00010110"; z_correct<="1111011100010000";
        when 6295 => y_in <= "10011000"; x_in <= "00010111"; z_correct<="1111011010101000";
        when 6296 => y_in <= "10011000"; x_in <= "00011000"; z_correct<="1111011001000000";
        when 6297 => y_in <= "10011000"; x_in <= "00011001"; z_correct<="1111010111011000";
        when 6298 => y_in <= "10011000"; x_in <= "00011010"; z_correct<="1111010101110000";
        when 6299 => y_in <= "10011000"; x_in <= "00011011"; z_correct<="1111010100001000";
        when 6300 => y_in <= "10011000"; x_in <= "00011100"; z_correct<="1111010010100000";
        when 6301 => y_in <= "10011000"; x_in <= "00011101"; z_correct<="1111010000111000";
        when 6302 => y_in <= "10011000"; x_in <= "00011110"; z_correct<="1111001111010000";
        when 6303 => y_in <= "10011000"; x_in <= "00011111"; z_correct<="1111001101101000";
        when 6304 => y_in <= "10011000"; x_in <= "00100000"; z_correct<="1111001100000000";
        when 6305 => y_in <= "10011000"; x_in <= "00100001"; z_correct<="1111001010011000";
        when 6306 => y_in <= "10011000"; x_in <= "00100010"; z_correct<="1111001000110000";
        when 6307 => y_in <= "10011000"; x_in <= "00100011"; z_correct<="1111000111001000";
        when 6308 => y_in <= "10011000"; x_in <= "00100100"; z_correct<="1111000101100000";
        when 6309 => y_in <= "10011000"; x_in <= "00100101"; z_correct<="1111000011111000";
        when 6310 => y_in <= "10011000"; x_in <= "00100110"; z_correct<="1111000010010000";
        when 6311 => y_in <= "10011000"; x_in <= "00100111"; z_correct<="1111000000101000";
        when 6312 => y_in <= "10011000"; x_in <= "00101000"; z_correct<="1110111111000000";
        when 6313 => y_in <= "10011000"; x_in <= "00101001"; z_correct<="1110111101011000";
        when 6314 => y_in <= "10011000"; x_in <= "00101010"; z_correct<="1110111011110000";
        when 6315 => y_in <= "10011000"; x_in <= "00101011"; z_correct<="1110111010001000";
        when 6316 => y_in <= "10011000"; x_in <= "00101100"; z_correct<="1110111000100000";
        when 6317 => y_in <= "10011000"; x_in <= "00101101"; z_correct<="1110110110111000";
        when 6318 => y_in <= "10011000"; x_in <= "00101110"; z_correct<="1110110101010000";
        when 6319 => y_in <= "10011000"; x_in <= "00101111"; z_correct<="1110110011101000";
        when 6320 => y_in <= "10011000"; x_in <= "00110000"; z_correct<="1110110010000000";
        when 6321 => y_in <= "10011000"; x_in <= "00110001"; z_correct<="1110110000011000";
        when 6322 => y_in <= "10011000"; x_in <= "00110010"; z_correct<="1110101110110000";
        when 6323 => y_in <= "10011000"; x_in <= "00110011"; z_correct<="1110101101001000";
        when 6324 => y_in <= "10011000"; x_in <= "00110100"; z_correct<="1110101011100000";
        when 6325 => y_in <= "10011000"; x_in <= "00110101"; z_correct<="1110101001111000";
        when 6326 => y_in <= "10011000"; x_in <= "00110110"; z_correct<="1110101000010000";
        when 6327 => y_in <= "10011000"; x_in <= "00110111"; z_correct<="1110100110101000";
        when 6328 => y_in <= "10011000"; x_in <= "00111000"; z_correct<="1110100101000000";
        when 6329 => y_in <= "10011000"; x_in <= "00111001"; z_correct<="1110100011011000";
        when 6330 => y_in <= "10011000"; x_in <= "00111010"; z_correct<="1110100001110000";
        when 6331 => y_in <= "10011000"; x_in <= "00111011"; z_correct<="1110100000001000";
        when 6332 => y_in <= "10011000"; x_in <= "00111100"; z_correct<="1110011110100000";
        when 6333 => y_in <= "10011000"; x_in <= "00111101"; z_correct<="1110011100111000";
        when 6334 => y_in <= "10011000"; x_in <= "00111110"; z_correct<="1110011011010000";
        when 6335 => y_in <= "10011000"; x_in <= "00111111"; z_correct<="1110011001101000";
        when 6336 => y_in <= "10011000"; x_in <= "01000000"; z_correct<="1110011000000000";
        when 6337 => y_in <= "10011000"; x_in <= "01000001"; z_correct<="1110010110011000";
        when 6338 => y_in <= "10011000"; x_in <= "01000010"; z_correct<="1110010100110000";
        when 6339 => y_in <= "10011000"; x_in <= "01000011"; z_correct<="1110010011001000";
        when 6340 => y_in <= "10011000"; x_in <= "01000100"; z_correct<="1110010001100000";
        when 6341 => y_in <= "10011000"; x_in <= "01000101"; z_correct<="1110001111111000";
        when 6342 => y_in <= "10011000"; x_in <= "01000110"; z_correct<="1110001110010000";
        when 6343 => y_in <= "10011000"; x_in <= "01000111"; z_correct<="1110001100101000";
        when 6344 => y_in <= "10011000"; x_in <= "01001000"; z_correct<="1110001011000000";
        when 6345 => y_in <= "10011000"; x_in <= "01001001"; z_correct<="1110001001011000";
        when 6346 => y_in <= "10011000"; x_in <= "01001010"; z_correct<="1110000111110000";
        when 6347 => y_in <= "10011000"; x_in <= "01001011"; z_correct<="1110000110001000";
        when 6348 => y_in <= "10011000"; x_in <= "01001100"; z_correct<="1110000100100000";
        when 6349 => y_in <= "10011000"; x_in <= "01001101"; z_correct<="1110000010111000";
        when 6350 => y_in <= "10011000"; x_in <= "01001110"; z_correct<="1110000001010000";
        when 6351 => y_in <= "10011000"; x_in <= "01001111"; z_correct<="1101111111101000";
        when 6352 => y_in <= "10011000"; x_in <= "01010000"; z_correct<="1101111110000000";
        when 6353 => y_in <= "10011000"; x_in <= "01010001"; z_correct<="1101111100011000";
        when 6354 => y_in <= "10011000"; x_in <= "01010010"; z_correct<="1101111010110000";
        when 6355 => y_in <= "10011000"; x_in <= "01010011"; z_correct<="1101111001001000";
        when 6356 => y_in <= "10011000"; x_in <= "01010100"; z_correct<="1101110111100000";
        when 6357 => y_in <= "10011000"; x_in <= "01010101"; z_correct<="1101110101111000";
        when 6358 => y_in <= "10011000"; x_in <= "01010110"; z_correct<="1101110100010000";
        when 6359 => y_in <= "10011000"; x_in <= "01010111"; z_correct<="1101110010101000";
        when 6360 => y_in <= "10011000"; x_in <= "01011000"; z_correct<="1101110001000000";
        when 6361 => y_in <= "10011000"; x_in <= "01011001"; z_correct<="1101101111011000";
        when 6362 => y_in <= "10011000"; x_in <= "01011010"; z_correct<="1101101101110000";
        when 6363 => y_in <= "10011000"; x_in <= "01011011"; z_correct<="1101101100001000";
        when 6364 => y_in <= "10011000"; x_in <= "01011100"; z_correct<="1101101010100000";
        when 6365 => y_in <= "10011000"; x_in <= "01011101"; z_correct<="1101101000111000";
        when 6366 => y_in <= "10011000"; x_in <= "01011110"; z_correct<="1101100111010000";
        when 6367 => y_in <= "10011000"; x_in <= "01011111"; z_correct<="1101100101101000";
        when 6368 => y_in <= "10011000"; x_in <= "01100000"; z_correct<="1101100100000000";
        when 6369 => y_in <= "10011000"; x_in <= "01100001"; z_correct<="1101100010011000";
        when 6370 => y_in <= "10011000"; x_in <= "01100010"; z_correct<="1101100000110000";
        when 6371 => y_in <= "10011000"; x_in <= "01100011"; z_correct<="1101011111001000";
        when 6372 => y_in <= "10011000"; x_in <= "01100100"; z_correct<="1101011101100000";
        when 6373 => y_in <= "10011000"; x_in <= "01100101"; z_correct<="1101011011111000";
        when 6374 => y_in <= "10011000"; x_in <= "01100110"; z_correct<="1101011010010000";
        when 6375 => y_in <= "10011000"; x_in <= "01100111"; z_correct<="1101011000101000";
        when 6376 => y_in <= "10011000"; x_in <= "01101000"; z_correct<="1101010111000000";
        when 6377 => y_in <= "10011000"; x_in <= "01101001"; z_correct<="1101010101011000";
        when 6378 => y_in <= "10011000"; x_in <= "01101010"; z_correct<="1101010011110000";
        when 6379 => y_in <= "10011000"; x_in <= "01101011"; z_correct<="1101010010001000";
        when 6380 => y_in <= "10011000"; x_in <= "01101100"; z_correct<="1101010000100000";
        when 6381 => y_in <= "10011000"; x_in <= "01101101"; z_correct<="1101001110111000";
        when 6382 => y_in <= "10011000"; x_in <= "01101110"; z_correct<="1101001101010000";
        when 6383 => y_in <= "10011000"; x_in <= "01101111"; z_correct<="1101001011101000";
        when 6384 => y_in <= "10011000"; x_in <= "01110000"; z_correct<="1101001010000000";
        when 6385 => y_in <= "10011000"; x_in <= "01110001"; z_correct<="1101001000011000";
        when 6386 => y_in <= "10011000"; x_in <= "01110010"; z_correct<="1101000110110000";
        when 6387 => y_in <= "10011000"; x_in <= "01110011"; z_correct<="1101000101001000";
        when 6388 => y_in <= "10011000"; x_in <= "01110100"; z_correct<="1101000011100000";
        when 6389 => y_in <= "10011000"; x_in <= "01110101"; z_correct<="1101000001111000";
        when 6390 => y_in <= "10011000"; x_in <= "01110110"; z_correct<="1101000000010000";
        when 6391 => y_in <= "10011000"; x_in <= "01110111"; z_correct<="1100111110101000";
        when 6392 => y_in <= "10011000"; x_in <= "01111000"; z_correct<="1100111101000000";
        when 6393 => y_in <= "10011000"; x_in <= "01111001"; z_correct<="1100111011011000";
        when 6394 => y_in <= "10011000"; x_in <= "01111010"; z_correct<="1100111001110000";
        when 6395 => y_in <= "10011000"; x_in <= "01111011"; z_correct<="1100111000001000";
        when 6396 => y_in <= "10011000"; x_in <= "01111100"; z_correct<="1100110110100000";
        when 6397 => y_in <= "10011000"; x_in <= "01111101"; z_correct<="1100110100111000";
        when 6398 => y_in <= "10011000"; x_in <= "01111110"; z_correct<="1100110011010000";
        when 6399 => y_in <= "10011000"; x_in <= "01111111"; z_correct<="1100110001101000";
        when 6400 => y_in <= "10011001"; x_in <= "10000000"; z_correct<="0011001110000000";
        when 6401 => y_in <= "10011001"; x_in <= "10000001"; z_correct<="0011001100011001";
        when 6402 => y_in <= "10011001"; x_in <= "10000010"; z_correct<="0011001010110010";
        when 6403 => y_in <= "10011001"; x_in <= "10000011"; z_correct<="0011001001001011";
        when 6404 => y_in <= "10011001"; x_in <= "10000100"; z_correct<="0011000111100100";
        when 6405 => y_in <= "10011001"; x_in <= "10000101"; z_correct<="0011000101111101";
        when 6406 => y_in <= "10011001"; x_in <= "10000110"; z_correct<="0011000100010110";
        when 6407 => y_in <= "10011001"; x_in <= "10000111"; z_correct<="0011000010101111";
        when 6408 => y_in <= "10011001"; x_in <= "10001000"; z_correct<="0011000001001000";
        when 6409 => y_in <= "10011001"; x_in <= "10001001"; z_correct<="0010111111100001";
        when 6410 => y_in <= "10011001"; x_in <= "10001010"; z_correct<="0010111101111010";
        when 6411 => y_in <= "10011001"; x_in <= "10001011"; z_correct<="0010111100010011";
        when 6412 => y_in <= "10011001"; x_in <= "10001100"; z_correct<="0010111010101100";
        when 6413 => y_in <= "10011001"; x_in <= "10001101"; z_correct<="0010111001000101";
        when 6414 => y_in <= "10011001"; x_in <= "10001110"; z_correct<="0010110111011110";
        when 6415 => y_in <= "10011001"; x_in <= "10001111"; z_correct<="0010110101110111";
        when 6416 => y_in <= "10011001"; x_in <= "10010000"; z_correct<="0010110100010000";
        when 6417 => y_in <= "10011001"; x_in <= "10010001"; z_correct<="0010110010101001";
        when 6418 => y_in <= "10011001"; x_in <= "10010010"; z_correct<="0010110001000010";
        when 6419 => y_in <= "10011001"; x_in <= "10010011"; z_correct<="0010101111011011";
        when 6420 => y_in <= "10011001"; x_in <= "10010100"; z_correct<="0010101101110100";
        when 6421 => y_in <= "10011001"; x_in <= "10010101"; z_correct<="0010101100001101";
        when 6422 => y_in <= "10011001"; x_in <= "10010110"; z_correct<="0010101010100110";
        when 6423 => y_in <= "10011001"; x_in <= "10010111"; z_correct<="0010101000111111";
        when 6424 => y_in <= "10011001"; x_in <= "10011000"; z_correct<="0010100111011000";
        when 6425 => y_in <= "10011001"; x_in <= "10011001"; z_correct<="0010100101110001";
        when 6426 => y_in <= "10011001"; x_in <= "10011010"; z_correct<="0010100100001010";
        when 6427 => y_in <= "10011001"; x_in <= "10011011"; z_correct<="0010100010100011";
        when 6428 => y_in <= "10011001"; x_in <= "10011100"; z_correct<="0010100000111100";
        when 6429 => y_in <= "10011001"; x_in <= "10011101"; z_correct<="0010011111010101";
        when 6430 => y_in <= "10011001"; x_in <= "10011110"; z_correct<="0010011101101110";
        when 6431 => y_in <= "10011001"; x_in <= "10011111"; z_correct<="0010011100000111";
        when 6432 => y_in <= "10011001"; x_in <= "10100000"; z_correct<="0010011010100000";
        when 6433 => y_in <= "10011001"; x_in <= "10100001"; z_correct<="0010011000111001";
        when 6434 => y_in <= "10011001"; x_in <= "10100010"; z_correct<="0010010111010010";
        when 6435 => y_in <= "10011001"; x_in <= "10100011"; z_correct<="0010010101101011";
        when 6436 => y_in <= "10011001"; x_in <= "10100100"; z_correct<="0010010100000100";
        when 6437 => y_in <= "10011001"; x_in <= "10100101"; z_correct<="0010010010011101";
        when 6438 => y_in <= "10011001"; x_in <= "10100110"; z_correct<="0010010000110110";
        when 6439 => y_in <= "10011001"; x_in <= "10100111"; z_correct<="0010001111001111";
        when 6440 => y_in <= "10011001"; x_in <= "10101000"; z_correct<="0010001101101000";
        when 6441 => y_in <= "10011001"; x_in <= "10101001"; z_correct<="0010001100000001";
        when 6442 => y_in <= "10011001"; x_in <= "10101010"; z_correct<="0010001010011010";
        when 6443 => y_in <= "10011001"; x_in <= "10101011"; z_correct<="0010001000110011";
        when 6444 => y_in <= "10011001"; x_in <= "10101100"; z_correct<="0010000111001100";
        when 6445 => y_in <= "10011001"; x_in <= "10101101"; z_correct<="0010000101100101";
        when 6446 => y_in <= "10011001"; x_in <= "10101110"; z_correct<="0010000011111110";
        when 6447 => y_in <= "10011001"; x_in <= "10101111"; z_correct<="0010000010010111";
        when 6448 => y_in <= "10011001"; x_in <= "10110000"; z_correct<="0010000000110000";
        when 6449 => y_in <= "10011001"; x_in <= "10110001"; z_correct<="0001111111001001";
        when 6450 => y_in <= "10011001"; x_in <= "10110010"; z_correct<="0001111101100010";
        when 6451 => y_in <= "10011001"; x_in <= "10110011"; z_correct<="0001111011111011";
        when 6452 => y_in <= "10011001"; x_in <= "10110100"; z_correct<="0001111010010100";
        when 6453 => y_in <= "10011001"; x_in <= "10110101"; z_correct<="0001111000101101";
        when 6454 => y_in <= "10011001"; x_in <= "10110110"; z_correct<="0001110111000110";
        when 6455 => y_in <= "10011001"; x_in <= "10110111"; z_correct<="0001110101011111";
        when 6456 => y_in <= "10011001"; x_in <= "10111000"; z_correct<="0001110011111000";
        when 6457 => y_in <= "10011001"; x_in <= "10111001"; z_correct<="0001110010010001";
        when 6458 => y_in <= "10011001"; x_in <= "10111010"; z_correct<="0001110000101010";
        when 6459 => y_in <= "10011001"; x_in <= "10111011"; z_correct<="0001101111000011";
        when 6460 => y_in <= "10011001"; x_in <= "10111100"; z_correct<="0001101101011100";
        when 6461 => y_in <= "10011001"; x_in <= "10111101"; z_correct<="0001101011110101";
        when 6462 => y_in <= "10011001"; x_in <= "10111110"; z_correct<="0001101010001110";
        when 6463 => y_in <= "10011001"; x_in <= "10111111"; z_correct<="0001101000100111";
        when 6464 => y_in <= "10011001"; x_in <= "11000000"; z_correct<="0001100111000000";
        when 6465 => y_in <= "10011001"; x_in <= "11000001"; z_correct<="0001100101011001";
        when 6466 => y_in <= "10011001"; x_in <= "11000010"; z_correct<="0001100011110010";
        when 6467 => y_in <= "10011001"; x_in <= "11000011"; z_correct<="0001100010001011";
        when 6468 => y_in <= "10011001"; x_in <= "11000100"; z_correct<="0001100000100100";
        when 6469 => y_in <= "10011001"; x_in <= "11000101"; z_correct<="0001011110111101";
        when 6470 => y_in <= "10011001"; x_in <= "11000110"; z_correct<="0001011101010110";
        when 6471 => y_in <= "10011001"; x_in <= "11000111"; z_correct<="0001011011101111";
        when 6472 => y_in <= "10011001"; x_in <= "11001000"; z_correct<="0001011010001000";
        when 6473 => y_in <= "10011001"; x_in <= "11001001"; z_correct<="0001011000100001";
        when 6474 => y_in <= "10011001"; x_in <= "11001010"; z_correct<="0001010110111010";
        when 6475 => y_in <= "10011001"; x_in <= "11001011"; z_correct<="0001010101010011";
        when 6476 => y_in <= "10011001"; x_in <= "11001100"; z_correct<="0001010011101100";
        when 6477 => y_in <= "10011001"; x_in <= "11001101"; z_correct<="0001010010000101";
        when 6478 => y_in <= "10011001"; x_in <= "11001110"; z_correct<="0001010000011110";
        when 6479 => y_in <= "10011001"; x_in <= "11001111"; z_correct<="0001001110110111";
        when 6480 => y_in <= "10011001"; x_in <= "11010000"; z_correct<="0001001101010000";
        when 6481 => y_in <= "10011001"; x_in <= "11010001"; z_correct<="0001001011101001";
        when 6482 => y_in <= "10011001"; x_in <= "11010010"; z_correct<="0001001010000010";
        when 6483 => y_in <= "10011001"; x_in <= "11010011"; z_correct<="0001001000011011";
        when 6484 => y_in <= "10011001"; x_in <= "11010100"; z_correct<="0001000110110100";
        when 6485 => y_in <= "10011001"; x_in <= "11010101"; z_correct<="0001000101001101";
        when 6486 => y_in <= "10011001"; x_in <= "11010110"; z_correct<="0001000011100110";
        when 6487 => y_in <= "10011001"; x_in <= "11010111"; z_correct<="0001000001111111";
        when 6488 => y_in <= "10011001"; x_in <= "11011000"; z_correct<="0001000000011000";
        when 6489 => y_in <= "10011001"; x_in <= "11011001"; z_correct<="0000111110110001";
        when 6490 => y_in <= "10011001"; x_in <= "11011010"; z_correct<="0000111101001010";
        when 6491 => y_in <= "10011001"; x_in <= "11011011"; z_correct<="0000111011100011";
        when 6492 => y_in <= "10011001"; x_in <= "11011100"; z_correct<="0000111001111100";
        when 6493 => y_in <= "10011001"; x_in <= "11011101"; z_correct<="0000111000010101";
        when 6494 => y_in <= "10011001"; x_in <= "11011110"; z_correct<="0000110110101110";
        when 6495 => y_in <= "10011001"; x_in <= "11011111"; z_correct<="0000110101000111";
        when 6496 => y_in <= "10011001"; x_in <= "11100000"; z_correct<="0000110011100000";
        when 6497 => y_in <= "10011001"; x_in <= "11100001"; z_correct<="0000110001111001";
        when 6498 => y_in <= "10011001"; x_in <= "11100010"; z_correct<="0000110000010010";
        when 6499 => y_in <= "10011001"; x_in <= "11100011"; z_correct<="0000101110101011";
        when 6500 => y_in <= "10011001"; x_in <= "11100100"; z_correct<="0000101101000100";
        when 6501 => y_in <= "10011001"; x_in <= "11100101"; z_correct<="0000101011011101";
        when 6502 => y_in <= "10011001"; x_in <= "11100110"; z_correct<="0000101001110110";
        when 6503 => y_in <= "10011001"; x_in <= "11100111"; z_correct<="0000101000001111";
        when 6504 => y_in <= "10011001"; x_in <= "11101000"; z_correct<="0000100110101000";
        when 6505 => y_in <= "10011001"; x_in <= "11101001"; z_correct<="0000100101000001";
        when 6506 => y_in <= "10011001"; x_in <= "11101010"; z_correct<="0000100011011010";
        when 6507 => y_in <= "10011001"; x_in <= "11101011"; z_correct<="0000100001110011";
        when 6508 => y_in <= "10011001"; x_in <= "11101100"; z_correct<="0000100000001100";
        when 6509 => y_in <= "10011001"; x_in <= "11101101"; z_correct<="0000011110100101";
        when 6510 => y_in <= "10011001"; x_in <= "11101110"; z_correct<="0000011100111110";
        when 6511 => y_in <= "10011001"; x_in <= "11101111"; z_correct<="0000011011010111";
        when 6512 => y_in <= "10011001"; x_in <= "11110000"; z_correct<="0000011001110000";
        when 6513 => y_in <= "10011001"; x_in <= "11110001"; z_correct<="0000011000001001";
        when 6514 => y_in <= "10011001"; x_in <= "11110010"; z_correct<="0000010110100010";
        when 6515 => y_in <= "10011001"; x_in <= "11110011"; z_correct<="0000010100111011";
        when 6516 => y_in <= "10011001"; x_in <= "11110100"; z_correct<="0000010011010100";
        when 6517 => y_in <= "10011001"; x_in <= "11110101"; z_correct<="0000010001101101";
        when 6518 => y_in <= "10011001"; x_in <= "11110110"; z_correct<="0000010000000110";
        when 6519 => y_in <= "10011001"; x_in <= "11110111"; z_correct<="0000001110011111";
        when 6520 => y_in <= "10011001"; x_in <= "11111000"; z_correct<="0000001100111000";
        when 6521 => y_in <= "10011001"; x_in <= "11111001"; z_correct<="0000001011010001";
        when 6522 => y_in <= "10011001"; x_in <= "11111010"; z_correct<="0000001001101010";
        when 6523 => y_in <= "10011001"; x_in <= "11111011"; z_correct<="0000001000000011";
        when 6524 => y_in <= "10011001"; x_in <= "11111100"; z_correct<="0000000110011100";
        when 6525 => y_in <= "10011001"; x_in <= "11111101"; z_correct<="0000000100110101";
        when 6526 => y_in <= "10011001"; x_in <= "11111110"; z_correct<="0000000011001110";
        when 6527 => y_in <= "10011001"; x_in <= "11111111"; z_correct<="0000000001100111";
        when 6528 => y_in <= "10011001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 6529 => y_in <= "10011001"; x_in <= "00000001"; z_correct<="1111111110011001";
        when 6530 => y_in <= "10011001"; x_in <= "00000010"; z_correct<="1111111100110010";
        when 6531 => y_in <= "10011001"; x_in <= "00000011"; z_correct<="1111111011001011";
        when 6532 => y_in <= "10011001"; x_in <= "00000100"; z_correct<="1111111001100100";
        when 6533 => y_in <= "10011001"; x_in <= "00000101"; z_correct<="1111110111111101";
        when 6534 => y_in <= "10011001"; x_in <= "00000110"; z_correct<="1111110110010110";
        when 6535 => y_in <= "10011001"; x_in <= "00000111"; z_correct<="1111110100101111";
        when 6536 => y_in <= "10011001"; x_in <= "00001000"; z_correct<="1111110011001000";
        when 6537 => y_in <= "10011001"; x_in <= "00001001"; z_correct<="1111110001100001";
        when 6538 => y_in <= "10011001"; x_in <= "00001010"; z_correct<="1111101111111010";
        when 6539 => y_in <= "10011001"; x_in <= "00001011"; z_correct<="1111101110010011";
        when 6540 => y_in <= "10011001"; x_in <= "00001100"; z_correct<="1111101100101100";
        when 6541 => y_in <= "10011001"; x_in <= "00001101"; z_correct<="1111101011000101";
        when 6542 => y_in <= "10011001"; x_in <= "00001110"; z_correct<="1111101001011110";
        when 6543 => y_in <= "10011001"; x_in <= "00001111"; z_correct<="1111100111110111";
        when 6544 => y_in <= "10011001"; x_in <= "00010000"; z_correct<="1111100110010000";
        when 6545 => y_in <= "10011001"; x_in <= "00010001"; z_correct<="1111100100101001";
        when 6546 => y_in <= "10011001"; x_in <= "00010010"; z_correct<="1111100011000010";
        when 6547 => y_in <= "10011001"; x_in <= "00010011"; z_correct<="1111100001011011";
        when 6548 => y_in <= "10011001"; x_in <= "00010100"; z_correct<="1111011111110100";
        when 6549 => y_in <= "10011001"; x_in <= "00010101"; z_correct<="1111011110001101";
        when 6550 => y_in <= "10011001"; x_in <= "00010110"; z_correct<="1111011100100110";
        when 6551 => y_in <= "10011001"; x_in <= "00010111"; z_correct<="1111011010111111";
        when 6552 => y_in <= "10011001"; x_in <= "00011000"; z_correct<="1111011001011000";
        when 6553 => y_in <= "10011001"; x_in <= "00011001"; z_correct<="1111010111110001";
        when 6554 => y_in <= "10011001"; x_in <= "00011010"; z_correct<="1111010110001010";
        when 6555 => y_in <= "10011001"; x_in <= "00011011"; z_correct<="1111010100100011";
        when 6556 => y_in <= "10011001"; x_in <= "00011100"; z_correct<="1111010010111100";
        when 6557 => y_in <= "10011001"; x_in <= "00011101"; z_correct<="1111010001010101";
        when 6558 => y_in <= "10011001"; x_in <= "00011110"; z_correct<="1111001111101110";
        when 6559 => y_in <= "10011001"; x_in <= "00011111"; z_correct<="1111001110000111";
        when 6560 => y_in <= "10011001"; x_in <= "00100000"; z_correct<="1111001100100000";
        when 6561 => y_in <= "10011001"; x_in <= "00100001"; z_correct<="1111001010111001";
        when 6562 => y_in <= "10011001"; x_in <= "00100010"; z_correct<="1111001001010010";
        when 6563 => y_in <= "10011001"; x_in <= "00100011"; z_correct<="1111000111101011";
        when 6564 => y_in <= "10011001"; x_in <= "00100100"; z_correct<="1111000110000100";
        when 6565 => y_in <= "10011001"; x_in <= "00100101"; z_correct<="1111000100011101";
        when 6566 => y_in <= "10011001"; x_in <= "00100110"; z_correct<="1111000010110110";
        when 6567 => y_in <= "10011001"; x_in <= "00100111"; z_correct<="1111000001001111";
        when 6568 => y_in <= "10011001"; x_in <= "00101000"; z_correct<="1110111111101000";
        when 6569 => y_in <= "10011001"; x_in <= "00101001"; z_correct<="1110111110000001";
        when 6570 => y_in <= "10011001"; x_in <= "00101010"; z_correct<="1110111100011010";
        when 6571 => y_in <= "10011001"; x_in <= "00101011"; z_correct<="1110111010110011";
        when 6572 => y_in <= "10011001"; x_in <= "00101100"; z_correct<="1110111001001100";
        when 6573 => y_in <= "10011001"; x_in <= "00101101"; z_correct<="1110110111100101";
        when 6574 => y_in <= "10011001"; x_in <= "00101110"; z_correct<="1110110101111110";
        when 6575 => y_in <= "10011001"; x_in <= "00101111"; z_correct<="1110110100010111";
        when 6576 => y_in <= "10011001"; x_in <= "00110000"; z_correct<="1110110010110000";
        when 6577 => y_in <= "10011001"; x_in <= "00110001"; z_correct<="1110110001001001";
        when 6578 => y_in <= "10011001"; x_in <= "00110010"; z_correct<="1110101111100010";
        when 6579 => y_in <= "10011001"; x_in <= "00110011"; z_correct<="1110101101111011";
        when 6580 => y_in <= "10011001"; x_in <= "00110100"; z_correct<="1110101100010100";
        when 6581 => y_in <= "10011001"; x_in <= "00110101"; z_correct<="1110101010101101";
        when 6582 => y_in <= "10011001"; x_in <= "00110110"; z_correct<="1110101001000110";
        when 6583 => y_in <= "10011001"; x_in <= "00110111"; z_correct<="1110100111011111";
        when 6584 => y_in <= "10011001"; x_in <= "00111000"; z_correct<="1110100101111000";
        when 6585 => y_in <= "10011001"; x_in <= "00111001"; z_correct<="1110100100010001";
        when 6586 => y_in <= "10011001"; x_in <= "00111010"; z_correct<="1110100010101010";
        when 6587 => y_in <= "10011001"; x_in <= "00111011"; z_correct<="1110100001000011";
        when 6588 => y_in <= "10011001"; x_in <= "00111100"; z_correct<="1110011111011100";
        when 6589 => y_in <= "10011001"; x_in <= "00111101"; z_correct<="1110011101110101";
        when 6590 => y_in <= "10011001"; x_in <= "00111110"; z_correct<="1110011100001110";
        when 6591 => y_in <= "10011001"; x_in <= "00111111"; z_correct<="1110011010100111";
        when 6592 => y_in <= "10011001"; x_in <= "01000000"; z_correct<="1110011001000000";
        when 6593 => y_in <= "10011001"; x_in <= "01000001"; z_correct<="1110010111011001";
        when 6594 => y_in <= "10011001"; x_in <= "01000010"; z_correct<="1110010101110010";
        when 6595 => y_in <= "10011001"; x_in <= "01000011"; z_correct<="1110010100001011";
        when 6596 => y_in <= "10011001"; x_in <= "01000100"; z_correct<="1110010010100100";
        when 6597 => y_in <= "10011001"; x_in <= "01000101"; z_correct<="1110010000111101";
        when 6598 => y_in <= "10011001"; x_in <= "01000110"; z_correct<="1110001111010110";
        when 6599 => y_in <= "10011001"; x_in <= "01000111"; z_correct<="1110001101101111";
        when 6600 => y_in <= "10011001"; x_in <= "01001000"; z_correct<="1110001100001000";
        when 6601 => y_in <= "10011001"; x_in <= "01001001"; z_correct<="1110001010100001";
        when 6602 => y_in <= "10011001"; x_in <= "01001010"; z_correct<="1110001000111010";
        when 6603 => y_in <= "10011001"; x_in <= "01001011"; z_correct<="1110000111010011";
        when 6604 => y_in <= "10011001"; x_in <= "01001100"; z_correct<="1110000101101100";
        when 6605 => y_in <= "10011001"; x_in <= "01001101"; z_correct<="1110000100000101";
        when 6606 => y_in <= "10011001"; x_in <= "01001110"; z_correct<="1110000010011110";
        when 6607 => y_in <= "10011001"; x_in <= "01001111"; z_correct<="1110000000110111";
        when 6608 => y_in <= "10011001"; x_in <= "01010000"; z_correct<="1101111111010000";
        when 6609 => y_in <= "10011001"; x_in <= "01010001"; z_correct<="1101111101101001";
        when 6610 => y_in <= "10011001"; x_in <= "01010010"; z_correct<="1101111100000010";
        when 6611 => y_in <= "10011001"; x_in <= "01010011"; z_correct<="1101111010011011";
        when 6612 => y_in <= "10011001"; x_in <= "01010100"; z_correct<="1101111000110100";
        when 6613 => y_in <= "10011001"; x_in <= "01010101"; z_correct<="1101110111001101";
        when 6614 => y_in <= "10011001"; x_in <= "01010110"; z_correct<="1101110101100110";
        when 6615 => y_in <= "10011001"; x_in <= "01010111"; z_correct<="1101110011111111";
        when 6616 => y_in <= "10011001"; x_in <= "01011000"; z_correct<="1101110010011000";
        when 6617 => y_in <= "10011001"; x_in <= "01011001"; z_correct<="1101110000110001";
        when 6618 => y_in <= "10011001"; x_in <= "01011010"; z_correct<="1101101111001010";
        when 6619 => y_in <= "10011001"; x_in <= "01011011"; z_correct<="1101101101100011";
        when 6620 => y_in <= "10011001"; x_in <= "01011100"; z_correct<="1101101011111100";
        when 6621 => y_in <= "10011001"; x_in <= "01011101"; z_correct<="1101101010010101";
        when 6622 => y_in <= "10011001"; x_in <= "01011110"; z_correct<="1101101000101110";
        when 6623 => y_in <= "10011001"; x_in <= "01011111"; z_correct<="1101100111000111";
        when 6624 => y_in <= "10011001"; x_in <= "01100000"; z_correct<="1101100101100000";
        when 6625 => y_in <= "10011001"; x_in <= "01100001"; z_correct<="1101100011111001";
        when 6626 => y_in <= "10011001"; x_in <= "01100010"; z_correct<="1101100010010010";
        when 6627 => y_in <= "10011001"; x_in <= "01100011"; z_correct<="1101100000101011";
        when 6628 => y_in <= "10011001"; x_in <= "01100100"; z_correct<="1101011111000100";
        when 6629 => y_in <= "10011001"; x_in <= "01100101"; z_correct<="1101011101011101";
        when 6630 => y_in <= "10011001"; x_in <= "01100110"; z_correct<="1101011011110110";
        when 6631 => y_in <= "10011001"; x_in <= "01100111"; z_correct<="1101011010001111";
        when 6632 => y_in <= "10011001"; x_in <= "01101000"; z_correct<="1101011000101000";
        when 6633 => y_in <= "10011001"; x_in <= "01101001"; z_correct<="1101010111000001";
        when 6634 => y_in <= "10011001"; x_in <= "01101010"; z_correct<="1101010101011010";
        when 6635 => y_in <= "10011001"; x_in <= "01101011"; z_correct<="1101010011110011";
        when 6636 => y_in <= "10011001"; x_in <= "01101100"; z_correct<="1101010010001100";
        when 6637 => y_in <= "10011001"; x_in <= "01101101"; z_correct<="1101010000100101";
        when 6638 => y_in <= "10011001"; x_in <= "01101110"; z_correct<="1101001110111110";
        when 6639 => y_in <= "10011001"; x_in <= "01101111"; z_correct<="1101001101010111";
        when 6640 => y_in <= "10011001"; x_in <= "01110000"; z_correct<="1101001011110000";
        when 6641 => y_in <= "10011001"; x_in <= "01110001"; z_correct<="1101001010001001";
        when 6642 => y_in <= "10011001"; x_in <= "01110010"; z_correct<="1101001000100010";
        when 6643 => y_in <= "10011001"; x_in <= "01110011"; z_correct<="1101000110111011";
        when 6644 => y_in <= "10011001"; x_in <= "01110100"; z_correct<="1101000101010100";
        when 6645 => y_in <= "10011001"; x_in <= "01110101"; z_correct<="1101000011101101";
        when 6646 => y_in <= "10011001"; x_in <= "01110110"; z_correct<="1101000010000110";
        when 6647 => y_in <= "10011001"; x_in <= "01110111"; z_correct<="1101000000011111";
        when 6648 => y_in <= "10011001"; x_in <= "01111000"; z_correct<="1100111110111000";
        when 6649 => y_in <= "10011001"; x_in <= "01111001"; z_correct<="1100111101010001";
        when 6650 => y_in <= "10011001"; x_in <= "01111010"; z_correct<="1100111011101010";
        when 6651 => y_in <= "10011001"; x_in <= "01111011"; z_correct<="1100111010000011";
        when 6652 => y_in <= "10011001"; x_in <= "01111100"; z_correct<="1100111000011100";
        when 6653 => y_in <= "10011001"; x_in <= "01111101"; z_correct<="1100110110110101";
        when 6654 => y_in <= "10011001"; x_in <= "01111110"; z_correct<="1100110101001110";
        when 6655 => y_in <= "10011001"; x_in <= "01111111"; z_correct<="1100110011100111";
        when 6656 => y_in <= "10011010"; x_in <= "10000000"; z_correct<="0011001100000000";
        when 6657 => y_in <= "10011010"; x_in <= "10000001"; z_correct<="0011001010011010";
        when 6658 => y_in <= "10011010"; x_in <= "10000010"; z_correct<="0011001000110100";
        when 6659 => y_in <= "10011010"; x_in <= "10000011"; z_correct<="0011000111001110";
        when 6660 => y_in <= "10011010"; x_in <= "10000100"; z_correct<="0011000101101000";
        when 6661 => y_in <= "10011010"; x_in <= "10000101"; z_correct<="0011000100000010";
        when 6662 => y_in <= "10011010"; x_in <= "10000110"; z_correct<="0011000010011100";
        when 6663 => y_in <= "10011010"; x_in <= "10000111"; z_correct<="0011000000110110";
        when 6664 => y_in <= "10011010"; x_in <= "10001000"; z_correct<="0010111111010000";
        when 6665 => y_in <= "10011010"; x_in <= "10001001"; z_correct<="0010111101101010";
        when 6666 => y_in <= "10011010"; x_in <= "10001010"; z_correct<="0010111100000100";
        when 6667 => y_in <= "10011010"; x_in <= "10001011"; z_correct<="0010111010011110";
        when 6668 => y_in <= "10011010"; x_in <= "10001100"; z_correct<="0010111000111000";
        when 6669 => y_in <= "10011010"; x_in <= "10001101"; z_correct<="0010110111010010";
        when 6670 => y_in <= "10011010"; x_in <= "10001110"; z_correct<="0010110101101100";
        when 6671 => y_in <= "10011010"; x_in <= "10001111"; z_correct<="0010110100000110";
        when 6672 => y_in <= "10011010"; x_in <= "10010000"; z_correct<="0010110010100000";
        when 6673 => y_in <= "10011010"; x_in <= "10010001"; z_correct<="0010110000111010";
        when 6674 => y_in <= "10011010"; x_in <= "10010010"; z_correct<="0010101111010100";
        when 6675 => y_in <= "10011010"; x_in <= "10010011"; z_correct<="0010101101101110";
        when 6676 => y_in <= "10011010"; x_in <= "10010100"; z_correct<="0010101100001000";
        when 6677 => y_in <= "10011010"; x_in <= "10010101"; z_correct<="0010101010100010";
        when 6678 => y_in <= "10011010"; x_in <= "10010110"; z_correct<="0010101000111100";
        when 6679 => y_in <= "10011010"; x_in <= "10010111"; z_correct<="0010100111010110";
        when 6680 => y_in <= "10011010"; x_in <= "10011000"; z_correct<="0010100101110000";
        when 6681 => y_in <= "10011010"; x_in <= "10011001"; z_correct<="0010100100001010";
        when 6682 => y_in <= "10011010"; x_in <= "10011010"; z_correct<="0010100010100100";
        when 6683 => y_in <= "10011010"; x_in <= "10011011"; z_correct<="0010100000111110";
        when 6684 => y_in <= "10011010"; x_in <= "10011100"; z_correct<="0010011111011000";
        when 6685 => y_in <= "10011010"; x_in <= "10011101"; z_correct<="0010011101110010";
        when 6686 => y_in <= "10011010"; x_in <= "10011110"; z_correct<="0010011100001100";
        when 6687 => y_in <= "10011010"; x_in <= "10011111"; z_correct<="0010011010100110";
        when 6688 => y_in <= "10011010"; x_in <= "10100000"; z_correct<="0010011001000000";
        when 6689 => y_in <= "10011010"; x_in <= "10100001"; z_correct<="0010010111011010";
        when 6690 => y_in <= "10011010"; x_in <= "10100010"; z_correct<="0010010101110100";
        when 6691 => y_in <= "10011010"; x_in <= "10100011"; z_correct<="0010010100001110";
        when 6692 => y_in <= "10011010"; x_in <= "10100100"; z_correct<="0010010010101000";
        when 6693 => y_in <= "10011010"; x_in <= "10100101"; z_correct<="0010010001000010";
        when 6694 => y_in <= "10011010"; x_in <= "10100110"; z_correct<="0010001111011100";
        when 6695 => y_in <= "10011010"; x_in <= "10100111"; z_correct<="0010001101110110";
        when 6696 => y_in <= "10011010"; x_in <= "10101000"; z_correct<="0010001100010000";
        when 6697 => y_in <= "10011010"; x_in <= "10101001"; z_correct<="0010001010101010";
        when 6698 => y_in <= "10011010"; x_in <= "10101010"; z_correct<="0010001001000100";
        when 6699 => y_in <= "10011010"; x_in <= "10101011"; z_correct<="0010000111011110";
        when 6700 => y_in <= "10011010"; x_in <= "10101100"; z_correct<="0010000101111000";
        when 6701 => y_in <= "10011010"; x_in <= "10101101"; z_correct<="0010000100010010";
        when 6702 => y_in <= "10011010"; x_in <= "10101110"; z_correct<="0010000010101100";
        when 6703 => y_in <= "10011010"; x_in <= "10101111"; z_correct<="0010000001000110";
        when 6704 => y_in <= "10011010"; x_in <= "10110000"; z_correct<="0001111111100000";
        when 6705 => y_in <= "10011010"; x_in <= "10110001"; z_correct<="0001111101111010";
        when 6706 => y_in <= "10011010"; x_in <= "10110010"; z_correct<="0001111100010100";
        when 6707 => y_in <= "10011010"; x_in <= "10110011"; z_correct<="0001111010101110";
        when 6708 => y_in <= "10011010"; x_in <= "10110100"; z_correct<="0001111001001000";
        when 6709 => y_in <= "10011010"; x_in <= "10110101"; z_correct<="0001110111100010";
        when 6710 => y_in <= "10011010"; x_in <= "10110110"; z_correct<="0001110101111100";
        when 6711 => y_in <= "10011010"; x_in <= "10110111"; z_correct<="0001110100010110";
        when 6712 => y_in <= "10011010"; x_in <= "10111000"; z_correct<="0001110010110000";
        when 6713 => y_in <= "10011010"; x_in <= "10111001"; z_correct<="0001110001001010";
        when 6714 => y_in <= "10011010"; x_in <= "10111010"; z_correct<="0001101111100100";
        when 6715 => y_in <= "10011010"; x_in <= "10111011"; z_correct<="0001101101111110";
        when 6716 => y_in <= "10011010"; x_in <= "10111100"; z_correct<="0001101100011000";
        when 6717 => y_in <= "10011010"; x_in <= "10111101"; z_correct<="0001101010110010";
        when 6718 => y_in <= "10011010"; x_in <= "10111110"; z_correct<="0001101001001100";
        when 6719 => y_in <= "10011010"; x_in <= "10111111"; z_correct<="0001100111100110";
        when 6720 => y_in <= "10011010"; x_in <= "11000000"; z_correct<="0001100110000000";
        when 6721 => y_in <= "10011010"; x_in <= "11000001"; z_correct<="0001100100011010";
        when 6722 => y_in <= "10011010"; x_in <= "11000010"; z_correct<="0001100010110100";
        when 6723 => y_in <= "10011010"; x_in <= "11000011"; z_correct<="0001100001001110";
        when 6724 => y_in <= "10011010"; x_in <= "11000100"; z_correct<="0001011111101000";
        when 6725 => y_in <= "10011010"; x_in <= "11000101"; z_correct<="0001011110000010";
        when 6726 => y_in <= "10011010"; x_in <= "11000110"; z_correct<="0001011100011100";
        when 6727 => y_in <= "10011010"; x_in <= "11000111"; z_correct<="0001011010110110";
        when 6728 => y_in <= "10011010"; x_in <= "11001000"; z_correct<="0001011001010000";
        when 6729 => y_in <= "10011010"; x_in <= "11001001"; z_correct<="0001010111101010";
        when 6730 => y_in <= "10011010"; x_in <= "11001010"; z_correct<="0001010110000100";
        when 6731 => y_in <= "10011010"; x_in <= "11001011"; z_correct<="0001010100011110";
        when 6732 => y_in <= "10011010"; x_in <= "11001100"; z_correct<="0001010010111000";
        when 6733 => y_in <= "10011010"; x_in <= "11001101"; z_correct<="0001010001010010";
        when 6734 => y_in <= "10011010"; x_in <= "11001110"; z_correct<="0001001111101100";
        when 6735 => y_in <= "10011010"; x_in <= "11001111"; z_correct<="0001001110000110";
        when 6736 => y_in <= "10011010"; x_in <= "11010000"; z_correct<="0001001100100000";
        when 6737 => y_in <= "10011010"; x_in <= "11010001"; z_correct<="0001001010111010";
        when 6738 => y_in <= "10011010"; x_in <= "11010010"; z_correct<="0001001001010100";
        when 6739 => y_in <= "10011010"; x_in <= "11010011"; z_correct<="0001000111101110";
        when 6740 => y_in <= "10011010"; x_in <= "11010100"; z_correct<="0001000110001000";
        when 6741 => y_in <= "10011010"; x_in <= "11010101"; z_correct<="0001000100100010";
        when 6742 => y_in <= "10011010"; x_in <= "11010110"; z_correct<="0001000010111100";
        when 6743 => y_in <= "10011010"; x_in <= "11010111"; z_correct<="0001000001010110";
        when 6744 => y_in <= "10011010"; x_in <= "11011000"; z_correct<="0000111111110000";
        when 6745 => y_in <= "10011010"; x_in <= "11011001"; z_correct<="0000111110001010";
        when 6746 => y_in <= "10011010"; x_in <= "11011010"; z_correct<="0000111100100100";
        when 6747 => y_in <= "10011010"; x_in <= "11011011"; z_correct<="0000111010111110";
        when 6748 => y_in <= "10011010"; x_in <= "11011100"; z_correct<="0000111001011000";
        when 6749 => y_in <= "10011010"; x_in <= "11011101"; z_correct<="0000110111110010";
        when 6750 => y_in <= "10011010"; x_in <= "11011110"; z_correct<="0000110110001100";
        when 6751 => y_in <= "10011010"; x_in <= "11011111"; z_correct<="0000110100100110";
        when 6752 => y_in <= "10011010"; x_in <= "11100000"; z_correct<="0000110011000000";
        when 6753 => y_in <= "10011010"; x_in <= "11100001"; z_correct<="0000110001011010";
        when 6754 => y_in <= "10011010"; x_in <= "11100010"; z_correct<="0000101111110100";
        when 6755 => y_in <= "10011010"; x_in <= "11100011"; z_correct<="0000101110001110";
        when 6756 => y_in <= "10011010"; x_in <= "11100100"; z_correct<="0000101100101000";
        when 6757 => y_in <= "10011010"; x_in <= "11100101"; z_correct<="0000101011000010";
        when 6758 => y_in <= "10011010"; x_in <= "11100110"; z_correct<="0000101001011100";
        when 6759 => y_in <= "10011010"; x_in <= "11100111"; z_correct<="0000100111110110";
        when 6760 => y_in <= "10011010"; x_in <= "11101000"; z_correct<="0000100110010000";
        when 6761 => y_in <= "10011010"; x_in <= "11101001"; z_correct<="0000100100101010";
        when 6762 => y_in <= "10011010"; x_in <= "11101010"; z_correct<="0000100011000100";
        when 6763 => y_in <= "10011010"; x_in <= "11101011"; z_correct<="0000100001011110";
        when 6764 => y_in <= "10011010"; x_in <= "11101100"; z_correct<="0000011111111000";
        when 6765 => y_in <= "10011010"; x_in <= "11101101"; z_correct<="0000011110010010";
        when 6766 => y_in <= "10011010"; x_in <= "11101110"; z_correct<="0000011100101100";
        when 6767 => y_in <= "10011010"; x_in <= "11101111"; z_correct<="0000011011000110";
        when 6768 => y_in <= "10011010"; x_in <= "11110000"; z_correct<="0000011001100000";
        when 6769 => y_in <= "10011010"; x_in <= "11110001"; z_correct<="0000010111111010";
        when 6770 => y_in <= "10011010"; x_in <= "11110010"; z_correct<="0000010110010100";
        when 6771 => y_in <= "10011010"; x_in <= "11110011"; z_correct<="0000010100101110";
        when 6772 => y_in <= "10011010"; x_in <= "11110100"; z_correct<="0000010011001000";
        when 6773 => y_in <= "10011010"; x_in <= "11110101"; z_correct<="0000010001100010";
        when 6774 => y_in <= "10011010"; x_in <= "11110110"; z_correct<="0000001111111100";
        when 6775 => y_in <= "10011010"; x_in <= "11110111"; z_correct<="0000001110010110";
        when 6776 => y_in <= "10011010"; x_in <= "11111000"; z_correct<="0000001100110000";
        when 6777 => y_in <= "10011010"; x_in <= "11111001"; z_correct<="0000001011001010";
        when 6778 => y_in <= "10011010"; x_in <= "11111010"; z_correct<="0000001001100100";
        when 6779 => y_in <= "10011010"; x_in <= "11111011"; z_correct<="0000000111111110";
        when 6780 => y_in <= "10011010"; x_in <= "11111100"; z_correct<="0000000110011000";
        when 6781 => y_in <= "10011010"; x_in <= "11111101"; z_correct<="0000000100110010";
        when 6782 => y_in <= "10011010"; x_in <= "11111110"; z_correct<="0000000011001100";
        when 6783 => y_in <= "10011010"; x_in <= "11111111"; z_correct<="0000000001100110";
        when 6784 => y_in <= "10011010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 6785 => y_in <= "10011010"; x_in <= "00000001"; z_correct<="1111111110011010";
        when 6786 => y_in <= "10011010"; x_in <= "00000010"; z_correct<="1111111100110100";
        when 6787 => y_in <= "10011010"; x_in <= "00000011"; z_correct<="1111111011001110";
        when 6788 => y_in <= "10011010"; x_in <= "00000100"; z_correct<="1111111001101000";
        when 6789 => y_in <= "10011010"; x_in <= "00000101"; z_correct<="1111111000000010";
        when 6790 => y_in <= "10011010"; x_in <= "00000110"; z_correct<="1111110110011100";
        when 6791 => y_in <= "10011010"; x_in <= "00000111"; z_correct<="1111110100110110";
        when 6792 => y_in <= "10011010"; x_in <= "00001000"; z_correct<="1111110011010000";
        when 6793 => y_in <= "10011010"; x_in <= "00001001"; z_correct<="1111110001101010";
        when 6794 => y_in <= "10011010"; x_in <= "00001010"; z_correct<="1111110000000100";
        when 6795 => y_in <= "10011010"; x_in <= "00001011"; z_correct<="1111101110011110";
        when 6796 => y_in <= "10011010"; x_in <= "00001100"; z_correct<="1111101100111000";
        when 6797 => y_in <= "10011010"; x_in <= "00001101"; z_correct<="1111101011010010";
        when 6798 => y_in <= "10011010"; x_in <= "00001110"; z_correct<="1111101001101100";
        when 6799 => y_in <= "10011010"; x_in <= "00001111"; z_correct<="1111101000000110";
        when 6800 => y_in <= "10011010"; x_in <= "00010000"; z_correct<="1111100110100000";
        when 6801 => y_in <= "10011010"; x_in <= "00010001"; z_correct<="1111100100111010";
        when 6802 => y_in <= "10011010"; x_in <= "00010010"; z_correct<="1111100011010100";
        when 6803 => y_in <= "10011010"; x_in <= "00010011"; z_correct<="1111100001101110";
        when 6804 => y_in <= "10011010"; x_in <= "00010100"; z_correct<="1111100000001000";
        when 6805 => y_in <= "10011010"; x_in <= "00010101"; z_correct<="1111011110100010";
        when 6806 => y_in <= "10011010"; x_in <= "00010110"; z_correct<="1111011100111100";
        when 6807 => y_in <= "10011010"; x_in <= "00010111"; z_correct<="1111011011010110";
        when 6808 => y_in <= "10011010"; x_in <= "00011000"; z_correct<="1111011001110000";
        when 6809 => y_in <= "10011010"; x_in <= "00011001"; z_correct<="1111011000001010";
        when 6810 => y_in <= "10011010"; x_in <= "00011010"; z_correct<="1111010110100100";
        when 6811 => y_in <= "10011010"; x_in <= "00011011"; z_correct<="1111010100111110";
        when 6812 => y_in <= "10011010"; x_in <= "00011100"; z_correct<="1111010011011000";
        when 6813 => y_in <= "10011010"; x_in <= "00011101"; z_correct<="1111010001110010";
        when 6814 => y_in <= "10011010"; x_in <= "00011110"; z_correct<="1111010000001100";
        when 6815 => y_in <= "10011010"; x_in <= "00011111"; z_correct<="1111001110100110";
        when 6816 => y_in <= "10011010"; x_in <= "00100000"; z_correct<="1111001101000000";
        when 6817 => y_in <= "10011010"; x_in <= "00100001"; z_correct<="1111001011011010";
        when 6818 => y_in <= "10011010"; x_in <= "00100010"; z_correct<="1111001001110100";
        when 6819 => y_in <= "10011010"; x_in <= "00100011"; z_correct<="1111001000001110";
        when 6820 => y_in <= "10011010"; x_in <= "00100100"; z_correct<="1111000110101000";
        when 6821 => y_in <= "10011010"; x_in <= "00100101"; z_correct<="1111000101000010";
        when 6822 => y_in <= "10011010"; x_in <= "00100110"; z_correct<="1111000011011100";
        when 6823 => y_in <= "10011010"; x_in <= "00100111"; z_correct<="1111000001110110";
        when 6824 => y_in <= "10011010"; x_in <= "00101000"; z_correct<="1111000000010000";
        when 6825 => y_in <= "10011010"; x_in <= "00101001"; z_correct<="1110111110101010";
        when 6826 => y_in <= "10011010"; x_in <= "00101010"; z_correct<="1110111101000100";
        when 6827 => y_in <= "10011010"; x_in <= "00101011"; z_correct<="1110111011011110";
        when 6828 => y_in <= "10011010"; x_in <= "00101100"; z_correct<="1110111001111000";
        when 6829 => y_in <= "10011010"; x_in <= "00101101"; z_correct<="1110111000010010";
        when 6830 => y_in <= "10011010"; x_in <= "00101110"; z_correct<="1110110110101100";
        when 6831 => y_in <= "10011010"; x_in <= "00101111"; z_correct<="1110110101000110";
        when 6832 => y_in <= "10011010"; x_in <= "00110000"; z_correct<="1110110011100000";
        when 6833 => y_in <= "10011010"; x_in <= "00110001"; z_correct<="1110110001111010";
        when 6834 => y_in <= "10011010"; x_in <= "00110010"; z_correct<="1110110000010100";
        when 6835 => y_in <= "10011010"; x_in <= "00110011"; z_correct<="1110101110101110";
        when 6836 => y_in <= "10011010"; x_in <= "00110100"; z_correct<="1110101101001000";
        when 6837 => y_in <= "10011010"; x_in <= "00110101"; z_correct<="1110101011100010";
        when 6838 => y_in <= "10011010"; x_in <= "00110110"; z_correct<="1110101001111100";
        when 6839 => y_in <= "10011010"; x_in <= "00110111"; z_correct<="1110101000010110";
        when 6840 => y_in <= "10011010"; x_in <= "00111000"; z_correct<="1110100110110000";
        when 6841 => y_in <= "10011010"; x_in <= "00111001"; z_correct<="1110100101001010";
        when 6842 => y_in <= "10011010"; x_in <= "00111010"; z_correct<="1110100011100100";
        when 6843 => y_in <= "10011010"; x_in <= "00111011"; z_correct<="1110100001111110";
        when 6844 => y_in <= "10011010"; x_in <= "00111100"; z_correct<="1110100000011000";
        when 6845 => y_in <= "10011010"; x_in <= "00111101"; z_correct<="1110011110110010";
        when 6846 => y_in <= "10011010"; x_in <= "00111110"; z_correct<="1110011101001100";
        when 6847 => y_in <= "10011010"; x_in <= "00111111"; z_correct<="1110011011100110";
        when 6848 => y_in <= "10011010"; x_in <= "01000000"; z_correct<="1110011010000000";
        when 6849 => y_in <= "10011010"; x_in <= "01000001"; z_correct<="1110011000011010";
        when 6850 => y_in <= "10011010"; x_in <= "01000010"; z_correct<="1110010110110100";
        when 6851 => y_in <= "10011010"; x_in <= "01000011"; z_correct<="1110010101001110";
        when 6852 => y_in <= "10011010"; x_in <= "01000100"; z_correct<="1110010011101000";
        when 6853 => y_in <= "10011010"; x_in <= "01000101"; z_correct<="1110010010000010";
        when 6854 => y_in <= "10011010"; x_in <= "01000110"; z_correct<="1110010000011100";
        when 6855 => y_in <= "10011010"; x_in <= "01000111"; z_correct<="1110001110110110";
        when 6856 => y_in <= "10011010"; x_in <= "01001000"; z_correct<="1110001101010000";
        when 6857 => y_in <= "10011010"; x_in <= "01001001"; z_correct<="1110001011101010";
        when 6858 => y_in <= "10011010"; x_in <= "01001010"; z_correct<="1110001010000100";
        when 6859 => y_in <= "10011010"; x_in <= "01001011"; z_correct<="1110001000011110";
        when 6860 => y_in <= "10011010"; x_in <= "01001100"; z_correct<="1110000110111000";
        when 6861 => y_in <= "10011010"; x_in <= "01001101"; z_correct<="1110000101010010";
        when 6862 => y_in <= "10011010"; x_in <= "01001110"; z_correct<="1110000011101100";
        when 6863 => y_in <= "10011010"; x_in <= "01001111"; z_correct<="1110000010000110";
        when 6864 => y_in <= "10011010"; x_in <= "01010000"; z_correct<="1110000000100000";
        when 6865 => y_in <= "10011010"; x_in <= "01010001"; z_correct<="1101111110111010";
        when 6866 => y_in <= "10011010"; x_in <= "01010010"; z_correct<="1101111101010100";
        when 6867 => y_in <= "10011010"; x_in <= "01010011"; z_correct<="1101111011101110";
        when 6868 => y_in <= "10011010"; x_in <= "01010100"; z_correct<="1101111010001000";
        when 6869 => y_in <= "10011010"; x_in <= "01010101"; z_correct<="1101111000100010";
        when 6870 => y_in <= "10011010"; x_in <= "01010110"; z_correct<="1101110110111100";
        when 6871 => y_in <= "10011010"; x_in <= "01010111"; z_correct<="1101110101010110";
        when 6872 => y_in <= "10011010"; x_in <= "01011000"; z_correct<="1101110011110000";
        when 6873 => y_in <= "10011010"; x_in <= "01011001"; z_correct<="1101110010001010";
        when 6874 => y_in <= "10011010"; x_in <= "01011010"; z_correct<="1101110000100100";
        when 6875 => y_in <= "10011010"; x_in <= "01011011"; z_correct<="1101101110111110";
        when 6876 => y_in <= "10011010"; x_in <= "01011100"; z_correct<="1101101101011000";
        when 6877 => y_in <= "10011010"; x_in <= "01011101"; z_correct<="1101101011110010";
        when 6878 => y_in <= "10011010"; x_in <= "01011110"; z_correct<="1101101010001100";
        when 6879 => y_in <= "10011010"; x_in <= "01011111"; z_correct<="1101101000100110";
        when 6880 => y_in <= "10011010"; x_in <= "01100000"; z_correct<="1101100111000000";
        when 6881 => y_in <= "10011010"; x_in <= "01100001"; z_correct<="1101100101011010";
        when 6882 => y_in <= "10011010"; x_in <= "01100010"; z_correct<="1101100011110100";
        when 6883 => y_in <= "10011010"; x_in <= "01100011"; z_correct<="1101100010001110";
        when 6884 => y_in <= "10011010"; x_in <= "01100100"; z_correct<="1101100000101000";
        when 6885 => y_in <= "10011010"; x_in <= "01100101"; z_correct<="1101011111000010";
        when 6886 => y_in <= "10011010"; x_in <= "01100110"; z_correct<="1101011101011100";
        when 6887 => y_in <= "10011010"; x_in <= "01100111"; z_correct<="1101011011110110";
        when 6888 => y_in <= "10011010"; x_in <= "01101000"; z_correct<="1101011010010000";
        when 6889 => y_in <= "10011010"; x_in <= "01101001"; z_correct<="1101011000101010";
        when 6890 => y_in <= "10011010"; x_in <= "01101010"; z_correct<="1101010111000100";
        when 6891 => y_in <= "10011010"; x_in <= "01101011"; z_correct<="1101010101011110";
        when 6892 => y_in <= "10011010"; x_in <= "01101100"; z_correct<="1101010011111000";
        when 6893 => y_in <= "10011010"; x_in <= "01101101"; z_correct<="1101010010010010";
        when 6894 => y_in <= "10011010"; x_in <= "01101110"; z_correct<="1101010000101100";
        when 6895 => y_in <= "10011010"; x_in <= "01101111"; z_correct<="1101001111000110";
        when 6896 => y_in <= "10011010"; x_in <= "01110000"; z_correct<="1101001101100000";
        when 6897 => y_in <= "10011010"; x_in <= "01110001"; z_correct<="1101001011111010";
        when 6898 => y_in <= "10011010"; x_in <= "01110010"; z_correct<="1101001010010100";
        when 6899 => y_in <= "10011010"; x_in <= "01110011"; z_correct<="1101001000101110";
        when 6900 => y_in <= "10011010"; x_in <= "01110100"; z_correct<="1101000111001000";
        when 6901 => y_in <= "10011010"; x_in <= "01110101"; z_correct<="1101000101100010";
        when 6902 => y_in <= "10011010"; x_in <= "01110110"; z_correct<="1101000011111100";
        when 6903 => y_in <= "10011010"; x_in <= "01110111"; z_correct<="1101000010010110";
        when 6904 => y_in <= "10011010"; x_in <= "01111000"; z_correct<="1101000000110000";
        when 6905 => y_in <= "10011010"; x_in <= "01111001"; z_correct<="1100111111001010";
        when 6906 => y_in <= "10011010"; x_in <= "01111010"; z_correct<="1100111101100100";
        when 6907 => y_in <= "10011010"; x_in <= "01111011"; z_correct<="1100111011111110";
        when 6908 => y_in <= "10011010"; x_in <= "01111100"; z_correct<="1100111010011000";
        when 6909 => y_in <= "10011010"; x_in <= "01111101"; z_correct<="1100111000110010";
        when 6910 => y_in <= "10011010"; x_in <= "01111110"; z_correct<="1100110111001100";
        when 6911 => y_in <= "10011010"; x_in <= "01111111"; z_correct<="1100110101100110";
        when 6912 => y_in <= "10011011"; x_in <= "10000000"; z_correct<="0011001010000000";
        when 6913 => y_in <= "10011011"; x_in <= "10000001"; z_correct<="0011001000011011";
        when 6914 => y_in <= "10011011"; x_in <= "10000010"; z_correct<="0011000110110110";
        when 6915 => y_in <= "10011011"; x_in <= "10000011"; z_correct<="0011000101010001";
        when 6916 => y_in <= "10011011"; x_in <= "10000100"; z_correct<="0011000011101100";
        when 6917 => y_in <= "10011011"; x_in <= "10000101"; z_correct<="0011000010000111";
        when 6918 => y_in <= "10011011"; x_in <= "10000110"; z_correct<="0011000000100010";
        when 6919 => y_in <= "10011011"; x_in <= "10000111"; z_correct<="0010111110111101";
        when 6920 => y_in <= "10011011"; x_in <= "10001000"; z_correct<="0010111101011000";
        when 6921 => y_in <= "10011011"; x_in <= "10001001"; z_correct<="0010111011110011";
        when 6922 => y_in <= "10011011"; x_in <= "10001010"; z_correct<="0010111010001110";
        when 6923 => y_in <= "10011011"; x_in <= "10001011"; z_correct<="0010111000101001";
        when 6924 => y_in <= "10011011"; x_in <= "10001100"; z_correct<="0010110111000100";
        when 6925 => y_in <= "10011011"; x_in <= "10001101"; z_correct<="0010110101011111";
        when 6926 => y_in <= "10011011"; x_in <= "10001110"; z_correct<="0010110011111010";
        when 6927 => y_in <= "10011011"; x_in <= "10001111"; z_correct<="0010110010010101";
        when 6928 => y_in <= "10011011"; x_in <= "10010000"; z_correct<="0010110000110000";
        when 6929 => y_in <= "10011011"; x_in <= "10010001"; z_correct<="0010101111001011";
        when 6930 => y_in <= "10011011"; x_in <= "10010010"; z_correct<="0010101101100110";
        when 6931 => y_in <= "10011011"; x_in <= "10010011"; z_correct<="0010101100000001";
        when 6932 => y_in <= "10011011"; x_in <= "10010100"; z_correct<="0010101010011100";
        when 6933 => y_in <= "10011011"; x_in <= "10010101"; z_correct<="0010101000110111";
        when 6934 => y_in <= "10011011"; x_in <= "10010110"; z_correct<="0010100111010010";
        when 6935 => y_in <= "10011011"; x_in <= "10010111"; z_correct<="0010100101101101";
        when 6936 => y_in <= "10011011"; x_in <= "10011000"; z_correct<="0010100100001000";
        when 6937 => y_in <= "10011011"; x_in <= "10011001"; z_correct<="0010100010100011";
        when 6938 => y_in <= "10011011"; x_in <= "10011010"; z_correct<="0010100000111110";
        when 6939 => y_in <= "10011011"; x_in <= "10011011"; z_correct<="0010011111011001";
        when 6940 => y_in <= "10011011"; x_in <= "10011100"; z_correct<="0010011101110100";
        when 6941 => y_in <= "10011011"; x_in <= "10011101"; z_correct<="0010011100001111";
        when 6942 => y_in <= "10011011"; x_in <= "10011110"; z_correct<="0010011010101010";
        when 6943 => y_in <= "10011011"; x_in <= "10011111"; z_correct<="0010011001000101";
        when 6944 => y_in <= "10011011"; x_in <= "10100000"; z_correct<="0010010111100000";
        when 6945 => y_in <= "10011011"; x_in <= "10100001"; z_correct<="0010010101111011";
        when 6946 => y_in <= "10011011"; x_in <= "10100010"; z_correct<="0010010100010110";
        when 6947 => y_in <= "10011011"; x_in <= "10100011"; z_correct<="0010010010110001";
        when 6948 => y_in <= "10011011"; x_in <= "10100100"; z_correct<="0010010001001100";
        when 6949 => y_in <= "10011011"; x_in <= "10100101"; z_correct<="0010001111100111";
        when 6950 => y_in <= "10011011"; x_in <= "10100110"; z_correct<="0010001110000010";
        when 6951 => y_in <= "10011011"; x_in <= "10100111"; z_correct<="0010001100011101";
        when 6952 => y_in <= "10011011"; x_in <= "10101000"; z_correct<="0010001010111000";
        when 6953 => y_in <= "10011011"; x_in <= "10101001"; z_correct<="0010001001010011";
        when 6954 => y_in <= "10011011"; x_in <= "10101010"; z_correct<="0010000111101110";
        when 6955 => y_in <= "10011011"; x_in <= "10101011"; z_correct<="0010000110001001";
        when 6956 => y_in <= "10011011"; x_in <= "10101100"; z_correct<="0010000100100100";
        when 6957 => y_in <= "10011011"; x_in <= "10101101"; z_correct<="0010000010111111";
        when 6958 => y_in <= "10011011"; x_in <= "10101110"; z_correct<="0010000001011010";
        when 6959 => y_in <= "10011011"; x_in <= "10101111"; z_correct<="0001111111110101";
        when 6960 => y_in <= "10011011"; x_in <= "10110000"; z_correct<="0001111110010000";
        when 6961 => y_in <= "10011011"; x_in <= "10110001"; z_correct<="0001111100101011";
        when 6962 => y_in <= "10011011"; x_in <= "10110010"; z_correct<="0001111011000110";
        when 6963 => y_in <= "10011011"; x_in <= "10110011"; z_correct<="0001111001100001";
        when 6964 => y_in <= "10011011"; x_in <= "10110100"; z_correct<="0001110111111100";
        when 6965 => y_in <= "10011011"; x_in <= "10110101"; z_correct<="0001110110010111";
        when 6966 => y_in <= "10011011"; x_in <= "10110110"; z_correct<="0001110100110010";
        when 6967 => y_in <= "10011011"; x_in <= "10110111"; z_correct<="0001110011001101";
        when 6968 => y_in <= "10011011"; x_in <= "10111000"; z_correct<="0001110001101000";
        when 6969 => y_in <= "10011011"; x_in <= "10111001"; z_correct<="0001110000000011";
        when 6970 => y_in <= "10011011"; x_in <= "10111010"; z_correct<="0001101110011110";
        when 6971 => y_in <= "10011011"; x_in <= "10111011"; z_correct<="0001101100111001";
        when 6972 => y_in <= "10011011"; x_in <= "10111100"; z_correct<="0001101011010100";
        when 6973 => y_in <= "10011011"; x_in <= "10111101"; z_correct<="0001101001101111";
        when 6974 => y_in <= "10011011"; x_in <= "10111110"; z_correct<="0001101000001010";
        when 6975 => y_in <= "10011011"; x_in <= "10111111"; z_correct<="0001100110100101";
        when 6976 => y_in <= "10011011"; x_in <= "11000000"; z_correct<="0001100101000000";
        when 6977 => y_in <= "10011011"; x_in <= "11000001"; z_correct<="0001100011011011";
        when 6978 => y_in <= "10011011"; x_in <= "11000010"; z_correct<="0001100001110110";
        when 6979 => y_in <= "10011011"; x_in <= "11000011"; z_correct<="0001100000010001";
        when 6980 => y_in <= "10011011"; x_in <= "11000100"; z_correct<="0001011110101100";
        when 6981 => y_in <= "10011011"; x_in <= "11000101"; z_correct<="0001011101000111";
        when 6982 => y_in <= "10011011"; x_in <= "11000110"; z_correct<="0001011011100010";
        when 6983 => y_in <= "10011011"; x_in <= "11000111"; z_correct<="0001011001111101";
        when 6984 => y_in <= "10011011"; x_in <= "11001000"; z_correct<="0001011000011000";
        when 6985 => y_in <= "10011011"; x_in <= "11001001"; z_correct<="0001010110110011";
        when 6986 => y_in <= "10011011"; x_in <= "11001010"; z_correct<="0001010101001110";
        when 6987 => y_in <= "10011011"; x_in <= "11001011"; z_correct<="0001010011101001";
        when 6988 => y_in <= "10011011"; x_in <= "11001100"; z_correct<="0001010010000100";
        when 6989 => y_in <= "10011011"; x_in <= "11001101"; z_correct<="0001010000011111";
        when 6990 => y_in <= "10011011"; x_in <= "11001110"; z_correct<="0001001110111010";
        when 6991 => y_in <= "10011011"; x_in <= "11001111"; z_correct<="0001001101010101";
        when 6992 => y_in <= "10011011"; x_in <= "11010000"; z_correct<="0001001011110000";
        when 6993 => y_in <= "10011011"; x_in <= "11010001"; z_correct<="0001001010001011";
        when 6994 => y_in <= "10011011"; x_in <= "11010010"; z_correct<="0001001000100110";
        when 6995 => y_in <= "10011011"; x_in <= "11010011"; z_correct<="0001000111000001";
        when 6996 => y_in <= "10011011"; x_in <= "11010100"; z_correct<="0001000101011100";
        when 6997 => y_in <= "10011011"; x_in <= "11010101"; z_correct<="0001000011110111";
        when 6998 => y_in <= "10011011"; x_in <= "11010110"; z_correct<="0001000010010010";
        when 6999 => y_in <= "10011011"; x_in <= "11010111"; z_correct<="0001000000101101";
        when 7000 => y_in <= "10011011"; x_in <= "11011000"; z_correct<="0000111111001000";
        when 7001 => y_in <= "10011011"; x_in <= "11011001"; z_correct<="0000111101100011";
        when 7002 => y_in <= "10011011"; x_in <= "11011010"; z_correct<="0000111011111110";
        when 7003 => y_in <= "10011011"; x_in <= "11011011"; z_correct<="0000111010011001";
        when 7004 => y_in <= "10011011"; x_in <= "11011100"; z_correct<="0000111000110100";
        when 7005 => y_in <= "10011011"; x_in <= "11011101"; z_correct<="0000110111001111";
        when 7006 => y_in <= "10011011"; x_in <= "11011110"; z_correct<="0000110101101010";
        when 7007 => y_in <= "10011011"; x_in <= "11011111"; z_correct<="0000110100000101";
        when 7008 => y_in <= "10011011"; x_in <= "11100000"; z_correct<="0000110010100000";
        when 7009 => y_in <= "10011011"; x_in <= "11100001"; z_correct<="0000110000111011";
        when 7010 => y_in <= "10011011"; x_in <= "11100010"; z_correct<="0000101111010110";
        when 7011 => y_in <= "10011011"; x_in <= "11100011"; z_correct<="0000101101110001";
        when 7012 => y_in <= "10011011"; x_in <= "11100100"; z_correct<="0000101100001100";
        when 7013 => y_in <= "10011011"; x_in <= "11100101"; z_correct<="0000101010100111";
        when 7014 => y_in <= "10011011"; x_in <= "11100110"; z_correct<="0000101001000010";
        when 7015 => y_in <= "10011011"; x_in <= "11100111"; z_correct<="0000100111011101";
        when 7016 => y_in <= "10011011"; x_in <= "11101000"; z_correct<="0000100101111000";
        when 7017 => y_in <= "10011011"; x_in <= "11101001"; z_correct<="0000100100010011";
        when 7018 => y_in <= "10011011"; x_in <= "11101010"; z_correct<="0000100010101110";
        when 7019 => y_in <= "10011011"; x_in <= "11101011"; z_correct<="0000100001001001";
        when 7020 => y_in <= "10011011"; x_in <= "11101100"; z_correct<="0000011111100100";
        when 7021 => y_in <= "10011011"; x_in <= "11101101"; z_correct<="0000011101111111";
        when 7022 => y_in <= "10011011"; x_in <= "11101110"; z_correct<="0000011100011010";
        when 7023 => y_in <= "10011011"; x_in <= "11101111"; z_correct<="0000011010110101";
        when 7024 => y_in <= "10011011"; x_in <= "11110000"; z_correct<="0000011001010000";
        when 7025 => y_in <= "10011011"; x_in <= "11110001"; z_correct<="0000010111101011";
        when 7026 => y_in <= "10011011"; x_in <= "11110010"; z_correct<="0000010110000110";
        when 7027 => y_in <= "10011011"; x_in <= "11110011"; z_correct<="0000010100100001";
        when 7028 => y_in <= "10011011"; x_in <= "11110100"; z_correct<="0000010010111100";
        when 7029 => y_in <= "10011011"; x_in <= "11110101"; z_correct<="0000010001010111";
        when 7030 => y_in <= "10011011"; x_in <= "11110110"; z_correct<="0000001111110010";
        when 7031 => y_in <= "10011011"; x_in <= "11110111"; z_correct<="0000001110001101";
        when 7032 => y_in <= "10011011"; x_in <= "11111000"; z_correct<="0000001100101000";
        when 7033 => y_in <= "10011011"; x_in <= "11111001"; z_correct<="0000001011000011";
        when 7034 => y_in <= "10011011"; x_in <= "11111010"; z_correct<="0000001001011110";
        when 7035 => y_in <= "10011011"; x_in <= "11111011"; z_correct<="0000000111111001";
        when 7036 => y_in <= "10011011"; x_in <= "11111100"; z_correct<="0000000110010100";
        when 7037 => y_in <= "10011011"; x_in <= "11111101"; z_correct<="0000000100101111";
        when 7038 => y_in <= "10011011"; x_in <= "11111110"; z_correct<="0000000011001010";
        when 7039 => y_in <= "10011011"; x_in <= "11111111"; z_correct<="0000000001100101";
        when 7040 => y_in <= "10011011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 7041 => y_in <= "10011011"; x_in <= "00000001"; z_correct<="1111111110011011";
        when 7042 => y_in <= "10011011"; x_in <= "00000010"; z_correct<="1111111100110110";
        when 7043 => y_in <= "10011011"; x_in <= "00000011"; z_correct<="1111111011010001";
        when 7044 => y_in <= "10011011"; x_in <= "00000100"; z_correct<="1111111001101100";
        when 7045 => y_in <= "10011011"; x_in <= "00000101"; z_correct<="1111111000000111";
        when 7046 => y_in <= "10011011"; x_in <= "00000110"; z_correct<="1111110110100010";
        when 7047 => y_in <= "10011011"; x_in <= "00000111"; z_correct<="1111110100111101";
        when 7048 => y_in <= "10011011"; x_in <= "00001000"; z_correct<="1111110011011000";
        when 7049 => y_in <= "10011011"; x_in <= "00001001"; z_correct<="1111110001110011";
        when 7050 => y_in <= "10011011"; x_in <= "00001010"; z_correct<="1111110000001110";
        when 7051 => y_in <= "10011011"; x_in <= "00001011"; z_correct<="1111101110101001";
        when 7052 => y_in <= "10011011"; x_in <= "00001100"; z_correct<="1111101101000100";
        when 7053 => y_in <= "10011011"; x_in <= "00001101"; z_correct<="1111101011011111";
        when 7054 => y_in <= "10011011"; x_in <= "00001110"; z_correct<="1111101001111010";
        when 7055 => y_in <= "10011011"; x_in <= "00001111"; z_correct<="1111101000010101";
        when 7056 => y_in <= "10011011"; x_in <= "00010000"; z_correct<="1111100110110000";
        when 7057 => y_in <= "10011011"; x_in <= "00010001"; z_correct<="1111100101001011";
        when 7058 => y_in <= "10011011"; x_in <= "00010010"; z_correct<="1111100011100110";
        when 7059 => y_in <= "10011011"; x_in <= "00010011"; z_correct<="1111100010000001";
        when 7060 => y_in <= "10011011"; x_in <= "00010100"; z_correct<="1111100000011100";
        when 7061 => y_in <= "10011011"; x_in <= "00010101"; z_correct<="1111011110110111";
        when 7062 => y_in <= "10011011"; x_in <= "00010110"; z_correct<="1111011101010010";
        when 7063 => y_in <= "10011011"; x_in <= "00010111"; z_correct<="1111011011101101";
        when 7064 => y_in <= "10011011"; x_in <= "00011000"; z_correct<="1111011010001000";
        when 7065 => y_in <= "10011011"; x_in <= "00011001"; z_correct<="1111011000100011";
        when 7066 => y_in <= "10011011"; x_in <= "00011010"; z_correct<="1111010110111110";
        when 7067 => y_in <= "10011011"; x_in <= "00011011"; z_correct<="1111010101011001";
        when 7068 => y_in <= "10011011"; x_in <= "00011100"; z_correct<="1111010011110100";
        when 7069 => y_in <= "10011011"; x_in <= "00011101"; z_correct<="1111010010001111";
        when 7070 => y_in <= "10011011"; x_in <= "00011110"; z_correct<="1111010000101010";
        when 7071 => y_in <= "10011011"; x_in <= "00011111"; z_correct<="1111001111000101";
        when 7072 => y_in <= "10011011"; x_in <= "00100000"; z_correct<="1111001101100000";
        when 7073 => y_in <= "10011011"; x_in <= "00100001"; z_correct<="1111001011111011";
        when 7074 => y_in <= "10011011"; x_in <= "00100010"; z_correct<="1111001010010110";
        when 7075 => y_in <= "10011011"; x_in <= "00100011"; z_correct<="1111001000110001";
        when 7076 => y_in <= "10011011"; x_in <= "00100100"; z_correct<="1111000111001100";
        when 7077 => y_in <= "10011011"; x_in <= "00100101"; z_correct<="1111000101100111";
        when 7078 => y_in <= "10011011"; x_in <= "00100110"; z_correct<="1111000100000010";
        when 7079 => y_in <= "10011011"; x_in <= "00100111"; z_correct<="1111000010011101";
        when 7080 => y_in <= "10011011"; x_in <= "00101000"; z_correct<="1111000000111000";
        when 7081 => y_in <= "10011011"; x_in <= "00101001"; z_correct<="1110111111010011";
        when 7082 => y_in <= "10011011"; x_in <= "00101010"; z_correct<="1110111101101110";
        when 7083 => y_in <= "10011011"; x_in <= "00101011"; z_correct<="1110111100001001";
        when 7084 => y_in <= "10011011"; x_in <= "00101100"; z_correct<="1110111010100100";
        when 7085 => y_in <= "10011011"; x_in <= "00101101"; z_correct<="1110111000111111";
        when 7086 => y_in <= "10011011"; x_in <= "00101110"; z_correct<="1110110111011010";
        when 7087 => y_in <= "10011011"; x_in <= "00101111"; z_correct<="1110110101110101";
        when 7088 => y_in <= "10011011"; x_in <= "00110000"; z_correct<="1110110100010000";
        when 7089 => y_in <= "10011011"; x_in <= "00110001"; z_correct<="1110110010101011";
        when 7090 => y_in <= "10011011"; x_in <= "00110010"; z_correct<="1110110001000110";
        when 7091 => y_in <= "10011011"; x_in <= "00110011"; z_correct<="1110101111100001";
        when 7092 => y_in <= "10011011"; x_in <= "00110100"; z_correct<="1110101101111100";
        when 7093 => y_in <= "10011011"; x_in <= "00110101"; z_correct<="1110101100010111";
        when 7094 => y_in <= "10011011"; x_in <= "00110110"; z_correct<="1110101010110010";
        when 7095 => y_in <= "10011011"; x_in <= "00110111"; z_correct<="1110101001001101";
        when 7096 => y_in <= "10011011"; x_in <= "00111000"; z_correct<="1110100111101000";
        when 7097 => y_in <= "10011011"; x_in <= "00111001"; z_correct<="1110100110000011";
        when 7098 => y_in <= "10011011"; x_in <= "00111010"; z_correct<="1110100100011110";
        when 7099 => y_in <= "10011011"; x_in <= "00111011"; z_correct<="1110100010111001";
        when 7100 => y_in <= "10011011"; x_in <= "00111100"; z_correct<="1110100001010100";
        when 7101 => y_in <= "10011011"; x_in <= "00111101"; z_correct<="1110011111101111";
        when 7102 => y_in <= "10011011"; x_in <= "00111110"; z_correct<="1110011110001010";
        when 7103 => y_in <= "10011011"; x_in <= "00111111"; z_correct<="1110011100100101";
        when 7104 => y_in <= "10011011"; x_in <= "01000000"; z_correct<="1110011011000000";
        when 7105 => y_in <= "10011011"; x_in <= "01000001"; z_correct<="1110011001011011";
        when 7106 => y_in <= "10011011"; x_in <= "01000010"; z_correct<="1110010111110110";
        when 7107 => y_in <= "10011011"; x_in <= "01000011"; z_correct<="1110010110010001";
        when 7108 => y_in <= "10011011"; x_in <= "01000100"; z_correct<="1110010100101100";
        when 7109 => y_in <= "10011011"; x_in <= "01000101"; z_correct<="1110010011000111";
        when 7110 => y_in <= "10011011"; x_in <= "01000110"; z_correct<="1110010001100010";
        when 7111 => y_in <= "10011011"; x_in <= "01000111"; z_correct<="1110001111111101";
        when 7112 => y_in <= "10011011"; x_in <= "01001000"; z_correct<="1110001110011000";
        when 7113 => y_in <= "10011011"; x_in <= "01001001"; z_correct<="1110001100110011";
        when 7114 => y_in <= "10011011"; x_in <= "01001010"; z_correct<="1110001011001110";
        when 7115 => y_in <= "10011011"; x_in <= "01001011"; z_correct<="1110001001101001";
        when 7116 => y_in <= "10011011"; x_in <= "01001100"; z_correct<="1110001000000100";
        when 7117 => y_in <= "10011011"; x_in <= "01001101"; z_correct<="1110000110011111";
        when 7118 => y_in <= "10011011"; x_in <= "01001110"; z_correct<="1110000100111010";
        when 7119 => y_in <= "10011011"; x_in <= "01001111"; z_correct<="1110000011010101";
        when 7120 => y_in <= "10011011"; x_in <= "01010000"; z_correct<="1110000001110000";
        when 7121 => y_in <= "10011011"; x_in <= "01010001"; z_correct<="1110000000001011";
        when 7122 => y_in <= "10011011"; x_in <= "01010010"; z_correct<="1101111110100110";
        when 7123 => y_in <= "10011011"; x_in <= "01010011"; z_correct<="1101111101000001";
        when 7124 => y_in <= "10011011"; x_in <= "01010100"; z_correct<="1101111011011100";
        when 7125 => y_in <= "10011011"; x_in <= "01010101"; z_correct<="1101111001110111";
        when 7126 => y_in <= "10011011"; x_in <= "01010110"; z_correct<="1101111000010010";
        when 7127 => y_in <= "10011011"; x_in <= "01010111"; z_correct<="1101110110101101";
        when 7128 => y_in <= "10011011"; x_in <= "01011000"; z_correct<="1101110101001000";
        when 7129 => y_in <= "10011011"; x_in <= "01011001"; z_correct<="1101110011100011";
        when 7130 => y_in <= "10011011"; x_in <= "01011010"; z_correct<="1101110001111110";
        when 7131 => y_in <= "10011011"; x_in <= "01011011"; z_correct<="1101110000011001";
        when 7132 => y_in <= "10011011"; x_in <= "01011100"; z_correct<="1101101110110100";
        when 7133 => y_in <= "10011011"; x_in <= "01011101"; z_correct<="1101101101001111";
        when 7134 => y_in <= "10011011"; x_in <= "01011110"; z_correct<="1101101011101010";
        when 7135 => y_in <= "10011011"; x_in <= "01011111"; z_correct<="1101101010000101";
        when 7136 => y_in <= "10011011"; x_in <= "01100000"; z_correct<="1101101000100000";
        when 7137 => y_in <= "10011011"; x_in <= "01100001"; z_correct<="1101100110111011";
        when 7138 => y_in <= "10011011"; x_in <= "01100010"; z_correct<="1101100101010110";
        when 7139 => y_in <= "10011011"; x_in <= "01100011"; z_correct<="1101100011110001";
        when 7140 => y_in <= "10011011"; x_in <= "01100100"; z_correct<="1101100010001100";
        when 7141 => y_in <= "10011011"; x_in <= "01100101"; z_correct<="1101100000100111";
        when 7142 => y_in <= "10011011"; x_in <= "01100110"; z_correct<="1101011111000010";
        when 7143 => y_in <= "10011011"; x_in <= "01100111"; z_correct<="1101011101011101";
        when 7144 => y_in <= "10011011"; x_in <= "01101000"; z_correct<="1101011011111000";
        when 7145 => y_in <= "10011011"; x_in <= "01101001"; z_correct<="1101011010010011";
        when 7146 => y_in <= "10011011"; x_in <= "01101010"; z_correct<="1101011000101110";
        when 7147 => y_in <= "10011011"; x_in <= "01101011"; z_correct<="1101010111001001";
        when 7148 => y_in <= "10011011"; x_in <= "01101100"; z_correct<="1101010101100100";
        when 7149 => y_in <= "10011011"; x_in <= "01101101"; z_correct<="1101010011111111";
        when 7150 => y_in <= "10011011"; x_in <= "01101110"; z_correct<="1101010010011010";
        when 7151 => y_in <= "10011011"; x_in <= "01101111"; z_correct<="1101010000110101";
        when 7152 => y_in <= "10011011"; x_in <= "01110000"; z_correct<="1101001111010000";
        when 7153 => y_in <= "10011011"; x_in <= "01110001"; z_correct<="1101001101101011";
        when 7154 => y_in <= "10011011"; x_in <= "01110010"; z_correct<="1101001100000110";
        when 7155 => y_in <= "10011011"; x_in <= "01110011"; z_correct<="1101001010100001";
        when 7156 => y_in <= "10011011"; x_in <= "01110100"; z_correct<="1101001000111100";
        when 7157 => y_in <= "10011011"; x_in <= "01110101"; z_correct<="1101000111010111";
        when 7158 => y_in <= "10011011"; x_in <= "01110110"; z_correct<="1101000101110010";
        when 7159 => y_in <= "10011011"; x_in <= "01110111"; z_correct<="1101000100001101";
        when 7160 => y_in <= "10011011"; x_in <= "01111000"; z_correct<="1101000010101000";
        when 7161 => y_in <= "10011011"; x_in <= "01111001"; z_correct<="1101000001000011";
        when 7162 => y_in <= "10011011"; x_in <= "01111010"; z_correct<="1100111111011110";
        when 7163 => y_in <= "10011011"; x_in <= "01111011"; z_correct<="1100111101111001";
        when 7164 => y_in <= "10011011"; x_in <= "01111100"; z_correct<="1100111100010100";
        when 7165 => y_in <= "10011011"; x_in <= "01111101"; z_correct<="1100111010101111";
        when 7166 => y_in <= "10011011"; x_in <= "01111110"; z_correct<="1100111001001010";
        when 7167 => y_in <= "10011011"; x_in <= "01111111"; z_correct<="1100110111100101";
        when 7168 => y_in <= "10011100"; x_in <= "10000000"; z_correct<="0011001000000000";
        when 7169 => y_in <= "10011100"; x_in <= "10000001"; z_correct<="0011000110011100";
        when 7170 => y_in <= "10011100"; x_in <= "10000010"; z_correct<="0011000100111000";
        when 7171 => y_in <= "10011100"; x_in <= "10000011"; z_correct<="0011000011010100";
        when 7172 => y_in <= "10011100"; x_in <= "10000100"; z_correct<="0011000001110000";
        when 7173 => y_in <= "10011100"; x_in <= "10000101"; z_correct<="0011000000001100";
        when 7174 => y_in <= "10011100"; x_in <= "10000110"; z_correct<="0010111110101000";
        when 7175 => y_in <= "10011100"; x_in <= "10000111"; z_correct<="0010111101000100";
        when 7176 => y_in <= "10011100"; x_in <= "10001000"; z_correct<="0010111011100000";
        when 7177 => y_in <= "10011100"; x_in <= "10001001"; z_correct<="0010111001111100";
        when 7178 => y_in <= "10011100"; x_in <= "10001010"; z_correct<="0010111000011000";
        when 7179 => y_in <= "10011100"; x_in <= "10001011"; z_correct<="0010110110110100";
        when 7180 => y_in <= "10011100"; x_in <= "10001100"; z_correct<="0010110101010000";
        when 7181 => y_in <= "10011100"; x_in <= "10001101"; z_correct<="0010110011101100";
        when 7182 => y_in <= "10011100"; x_in <= "10001110"; z_correct<="0010110010001000";
        when 7183 => y_in <= "10011100"; x_in <= "10001111"; z_correct<="0010110000100100";
        when 7184 => y_in <= "10011100"; x_in <= "10010000"; z_correct<="0010101111000000";
        when 7185 => y_in <= "10011100"; x_in <= "10010001"; z_correct<="0010101101011100";
        when 7186 => y_in <= "10011100"; x_in <= "10010010"; z_correct<="0010101011111000";
        when 7187 => y_in <= "10011100"; x_in <= "10010011"; z_correct<="0010101010010100";
        when 7188 => y_in <= "10011100"; x_in <= "10010100"; z_correct<="0010101000110000";
        when 7189 => y_in <= "10011100"; x_in <= "10010101"; z_correct<="0010100111001100";
        when 7190 => y_in <= "10011100"; x_in <= "10010110"; z_correct<="0010100101101000";
        when 7191 => y_in <= "10011100"; x_in <= "10010111"; z_correct<="0010100100000100";
        when 7192 => y_in <= "10011100"; x_in <= "10011000"; z_correct<="0010100010100000";
        when 7193 => y_in <= "10011100"; x_in <= "10011001"; z_correct<="0010100000111100";
        when 7194 => y_in <= "10011100"; x_in <= "10011010"; z_correct<="0010011111011000";
        when 7195 => y_in <= "10011100"; x_in <= "10011011"; z_correct<="0010011101110100";
        when 7196 => y_in <= "10011100"; x_in <= "10011100"; z_correct<="0010011100010000";
        when 7197 => y_in <= "10011100"; x_in <= "10011101"; z_correct<="0010011010101100";
        when 7198 => y_in <= "10011100"; x_in <= "10011110"; z_correct<="0010011001001000";
        when 7199 => y_in <= "10011100"; x_in <= "10011111"; z_correct<="0010010111100100";
        when 7200 => y_in <= "10011100"; x_in <= "10100000"; z_correct<="0010010110000000";
        when 7201 => y_in <= "10011100"; x_in <= "10100001"; z_correct<="0010010100011100";
        when 7202 => y_in <= "10011100"; x_in <= "10100010"; z_correct<="0010010010111000";
        when 7203 => y_in <= "10011100"; x_in <= "10100011"; z_correct<="0010010001010100";
        when 7204 => y_in <= "10011100"; x_in <= "10100100"; z_correct<="0010001111110000";
        when 7205 => y_in <= "10011100"; x_in <= "10100101"; z_correct<="0010001110001100";
        when 7206 => y_in <= "10011100"; x_in <= "10100110"; z_correct<="0010001100101000";
        when 7207 => y_in <= "10011100"; x_in <= "10100111"; z_correct<="0010001011000100";
        when 7208 => y_in <= "10011100"; x_in <= "10101000"; z_correct<="0010001001100000";
        when 7209 => y_in <= "10011100"; x_in <= "10101001"; z_correct<="0010000111111100";
        when 7210 => y_in <= "10011100"; x_in <= "10101010"; z_correct<="0010000110011000";
        when 7211 => y_in <= "10011100"; x_in <= "10101011"; z_correct<="0010000100110100";
        when 7212 => y_in <= "10011100"; x_in <= "10101100"; z_correct<="0010000011010000";
        when 7213 => y_in <= "10011100"; x_in <= "10101101"; z_correct<="0010000001101100";
        when 7214 => y_in <= "10011100"; x_in <= "10101110"; z_correct<="0010000000001000";
        when 7215 => y_in <= "10011100"; x_in <= "10101111"; z_correct<="0001111110100100";
        when 7216 => y_in <= "10011100"; x_in <= "10110000"; z_correct<="0001111101000000";
        when 7217 => y_in <= "10011100"; x_in <= "10110001"; z_correct<="0001111011011100";
        when 7218 => y_in <= "10011100"; x_in <= "10110010"; z_correct<="0001111001111000";
        when 7219 => y_in <= "10011100"; x_in <= "10110011"; z_correct<="0001111000010100";
        when 7220 => y_in <= "10011100"; x_in <= "10110100"; z_correct<="0001110110110000";
        when 7221 => y_in <= "10011100"; x_in <= "10110101"; z_correct<="0001110101001100";
        when 7222 => y_in <= "10011100"; x_in <= "10110110"; z_correct<="0001110011101000";
        when 7223 => y_in <= "10011100"; x_in <= "10110111"; z_correct<="0001110010000100";
        when 7224 => y_in <= "10011100"; x_in <= "10111000"; z_correct<="0001110000100000";
        when 7225 => y_in <= "10011100"; x_in <= "10111001"; z_correct<="0001101110111100";
        when 7226 => y_in <= "10011100"; x_in <= "10111010"; z_correct<="0001101101011000";
        when 7227 => y_in <= "10011100"; x_in <= "10111011"; z_correct<="0001101011110100";
        when 7228 => y_in <= "10011100"; x_in <= "10111100"; z_correct<="0001101010010000";
        when 7229 => y_in <= "10011100"; x_in <= "10111101"; z_correct<="0001101000101100";
        when 7230 => y_in <= "10011100"; x_in <= "10111110"; z_correct<="0001100111001000";
        when 7231 => y_in <= "10011100"; x_in <= "10111111"; z_correct<="0001100101100100";
        when 7232 => y_in <= "10011100"; x_in <= "11000000"; z_correct<="0001100100000000";
        when 7233 => y_in <= "10011100"; x_in <= "11000001"; z_correct<="0001100010011100";
        when 7234 => y_in <= "10011100"; x_in <= "11000010"; z_correct<="0001100000111000";
        when 7235 => y_in <= "10011100"; x_in <= "11000011"; z_correct<="0001011111010100";
        when 7236 => y_in <= "10011100"; x_in <= "11000100"; z_correct<="0001011101110000";
        when 7237 => y_in <= "10011100"; x_in <= "11000101"; z_correct<="0001011100001100";
        when 7238 => y_in <= "10011100"; x_in <= "11000110"; z_correct<="0001011010101000";
        when 7239 => y_in <= "10011100"; x_in <= "11000111"; z_correct<="0001011001000100";
        when 7240 => y_in <= "10011100"; x_in <= "11001000"; z_correct<="0001010111100000";
        when 7241 => y_in <= "10011100"; x_in <= "11001001"; z_correct<="0001010101111100";
        when 7242 => y_in <= "10011100"; x_in <= "11001010"; z_correct<="0001010100011000";
        when 7243 => y_in <= "10011100"; x_in <= "11001011"; z_correct<="0001010010110100";
        when 7244 => y_in <= "10011100"; x_in <= "11001100"; z_correct<="0001010001010000";
        when 7245 => y_in <= "10011100"; x_in <= "11001101"; z_correct<="0001001111101100";
        when 7246 => y_in <= "10011100"; x_in <= "11001110"; z_correct<="0001001110001000";
        when 7247 => y_in <= "10011100"; x_in <= "11001111"; z_correct<="0001001100100100";
        when 7248 => y_in <= "10011100"; x_in <= "11010000"; z_correct<="0001001011000000";
        when 7249 => y_in <= "10011100"; x_in <= "11010001"; z_correct<="0001001001011100";
        when 7250 => y_in <= "10011100"; x_in <= "11010010"; z_correct<="0001000111111000";
        when 7251 => y_in <= "10011100"; x_in <= "11010011"; z_correct<="0001000110010100";
        when 7252 => y_in <= "10011100"; x_in <= "11010100"; z_correct<="0001000100110000";
        when 7253 => y_in <= "10011100"; x_in <= "11010101"; z_correct<="0001000011001100";
        when 7254 => y_in <= "10011100"; x_in <= "11010110"; z_correct<="0001000001101000";
        when 7255 => y_in <= "10011100"; x_in <= "11010111"; z_correct<="0001000000000100";
        when 7256 => y_in <= "10011100"; x_in <= "11011000"; z_correct<="0000111110100000";
        when 7257 => y_in <= "10011100"; x_in <= "11011001"; z_correct<="0000111100111100";
        when 7258 => y_in <= "10011100"; x_in <= "11011010"; z_correct<="0000111011011000";
        when 7259 => y_in <= "10011100"; x_in <= "11011011"; z_correct<="0000111001110100";
        when 7260 => y_in <= "10011100"; x_in <= "11011100"; z_correct<="0000111000010000";
        when 7261 => y_in <= "10011100"; x_in <= "11011101"; z_correct<="0000110110101100";
        when 7262 => y_in <= "10011100"; x_in <= "11011110"; z_correct<="0000110101001000";
        when 7263 => y_in <= "10011100"; x_in <= "11011111"; z_correct<="0000110011100100";
        when 7264 => y_in <= "10011100"; x_in <= "11100000"; z_correct<="0000110010000000";
        when 7265 => y_in <= "10011100"; x_in <= "11100001"; z_correct<="0000110000011100";
        when 7266 => y_in <= "10011100"; x_in <= "11100010"; z_correct<="0000101110111000";
        when 7267 => y_in <= "10011100"; x_in <= "11100011"; z_correct<="0000101101010100";
        when 7268 => y_in <= "10011100"; x_in <= "11100100"; z_correct<="0000101011110000";
        when 7269 => y_in <= "10011100"; x_in <= "11100101"; z_correct<="0000101010001100";
        when 7270 => y_in <= "10011100"; x_in <= "11100110"; z_correct<="0000101000101000";
        when 7271 => y_in <= "10011100"; x_in <= "11100111"; z_correct<="0000100111000100";
        when 7272 => y_in <= "10011100"; x_in <= "11101000"; z_correct<="0000100101100000";
        when 7273 => y_in <= "10011100"; x_in <= "11101001"; z_correct<="0000100011111100";
        when 7274 => y_in <= "10011100"; x_in <= "11101010"; z_correct<="0000100010011000";
        when 7275 => y_in <= "10011100"; x_in <= "11101011"; z_correct<="0000100000110100";
        when 7276 => y_in <= "10011100"; x_in <= "11101100"; z_correct<="0000011111010000";
        when 7277 => y_in <= "10011100"; x_in <= "11101101"; z_correct<="0000011101101100";
        when 7278 => y_in <= "10011100"; x_in <= "11101110"; z_correct<="0000011100001000";
        when 7279 => y_in <= "10011100"; x_in <= "11101111"; z_correct<="0000011010100100";
        when 7280 => y_in <= "10011100"; x_in <= "11110000"; z_correct<="0000011001000000";
        when 7281 => y_in <= "10011100"; x_in <= "11110001"; z_correct<="0000010111011100";
        when 7282 => y_in <= "10011100"; x_in <= "11110010"; z_correct<="0000010101111000";
        when 7283 => y_in <= "10011100"; x_in <= "11110011"; z_correct<="0000010100010100";
        when 7284 => y_in <= "10011100"; x_in <= "11110100"; z_correct<="0000010010110000";
        when 7285 => y_in <= "10011100"; x_in <= "11110101"; z_correct<="0000010001001100";
        when 7286 => y_in <= "10011100"; x_in <= "11110110"; z_correct<="0000001111101000";
        when 7287 => y_in <= "10011100"; x_in <= "11110111"; z_correct<="0000001110000100";
        when 7288 => y_in <= "10011100"; x_in <= "11111000"; z_correct<="0000001100100000";
        when 7289 => y_in <= "10011100"; x_in <= "11111001"; z_correct<="0000001010111100";
        when 7290 => y_in <= "10011100"; x_in <= "11111010"; z_correct<="0000001001011000";
        when 7291 => y_in <= "10011100"; x_in <= "11111011"; z_correct<="0000000111110100";
        when 7292 => y_in <= "10011100"; x_in <= "11111100"; z_correct<="0000000110010000";
        when 7293 => y_in <= "10011100"; x_in <= "11111101"; z_correct<="0000000100101100";
        when 7294 => y_in <= "10011100"; x_in <= "11111110"; z_correct<="0000000011001000";
        when 7295 => y_in <= "10011100"; x_in <= "11111111"; z_correct<="0000000001100100";
        when 7296 => y_in <= "10011100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 7297 => y_in <= "10011100"; x_in <= "00000001"; z_correct<="1111111110011100";
        when 7298 => y_in <= "10011100"; x_in <= "00000010"; z_correct<="1111111100111000";
        when 7299 => y_in <= "10011100"; x_in <= "00000011"; z_correct<="1111111011010100";
        when 7300 => y_in <= "10011100"; x_in <= "00000100"; z_correct<="1111111001110000";
        when 7301 => y_in <= "10011100"; x_in <= "00000101"; z_correct<="1111111000001100";
        when 7302 => y_in <= "10011100"; x_in <= "00000110"; z_correct<="1111110110101000";
        when 7303 => y_in <= "10011100"; x_in <= "00000111"; z_correct<="1111110101000100";
        when 7304 => y_in <= "10011100"; x_in <= "00001000"; z_correct<="1111110011100000";
        when 7305 => y_in <= "10011100"; x_in <= "00001001"; z_correct<="1111110001111100";
        when 7306 => y_in <= "10011100"; x_in <= "00001010"; z_correct<="1111110000011000";
        when 7307 => y_in <= "10011100"; x_in <= "00001011"; z_correct<="1111101110110100";
        when 7308 => y_in <= "10011100"; x_in <= "00001100"; z_correct<="1111101101010000";
        when 7309 => y_in <= "10011100"; x_in <= "00001101"; z_correct<="1111101011101100";
        when 7310 => y_in <= "10011100"; x_in <= "00001110"; z_correct<="1111101010001000";
        when 7311 => y_in <= "10011100"; x_in <= "00001111"; z_correct<="1111101000100100";
        when 7312 => y_in <= "10011100"; x_in <= "00010000"; z_correct<="1111100111000000";
        when 7313 => y_in <= "10011100"; x_in <= "00010001"; z_correct<="1111100101011100";
        when 7314 => y_in <= "10011100"; x_in <= "00010010"; z_correct<="1111100011111000";
        when 7315 => y_in <= "10011100"; x_in <= "00010011"; z_correct<="1111100010010100";
        when 7316 => y_in <= "10011100"; x_in <= "00010100"; z_correct<="1111100000110000";
        when 7317 => y_in <= "10011100"; x_in <= "00010101"; z_correct<="1111011111001100";
        when 7318 => y_in <= "10011100"; x_in <= "00010110"; z_correct<="1111011101101000";
        when 7319 => y_in <= "10011100"; x_in <= "00010111"; z_correct<="1111011100000100";
        when 7320 => y_in <= "10011100"; x_in <= "00011000"; z_correct<="1111011010100000";
        when 7321 => y_in <= "10011100"; x_in <= "00011001"; z_correct<="1111011000111100";
        when 7322 => y_in <= "10011100"; x_in <= "00011010"; z_correct<="1111010111011000";
        when 7323 => y_in <= "10011100"; x_in <= "00011011"; z_correct<="1111010101110100";
        when 7324 => y_in <= "10011100"; x_in <= "00011100"; z_correct<="1111010100010000";
        when 7325 => y_in <= "10011100"; x_in <= "00011101"; z_correct<="1111010010101100";
        when 7326 => y_in <= "10011100"; x_in <= "00011110"; z_correct<="1111010001001000";
        when 7327 => y_in <= "10011100"; x_in <= "00011111"; z_correct<="1111001111100100";
        when 7328 => y_in <= "10011100"; x_in <= "00100000"; z_correct<="1111001110000000";
        when 7329 => y_in <= "10011100"; x_in <= "00100001"; z_correct<="1111001100011100";
        when 7330 => y_in <= "10011100"; x_in <= "00100010"; z_correct<="1111001010111000";
        when 7331 => y_in <= "10011100"; x_in <= "00100011"; z_correct<="1111001001010100";
        when 7332 => y_in <= "10011100"; x_in <= "00100100"; z_correct<="1111000111110000";
        when 7333 => y_in <= "10011100"; x_in <= "00100101"; z_correct<="1111000110001100";
        when 7334 => y_in <= "10011100"; x_in <= "00100110"; z_correct<="1111000100101000";
        when 7335 => y_in <= "10011100"; x_in <= "00100111"; z_correct<="1111000011000100";
        when 7336 => y_in <= "10011100"; x_in <= "00101000"; z_correct<="1111000001100000";
        when 7337 => y_in <= "10011100"; x_in <= "00101001"; z_correct<="1110111111111100";
        when 7338 => y_in <= "10011100"; x_in <= "00101010"; z_correct<="1110111110011000";
        when 7339 => y_in <= "10011100"; x_in <= "00101011"; z_correct<="1110111100110100";
        when 7340 => y_in <= "10011100"; x_in <= "00101100"; z_correct<="1110111011010000";
        when 7341 => y_in <= "10011100"; x_in <= "00101101"; z_correct<="1110111001101100";
        when 7342 => y_in <= "10011100"; x_in <= "00101110"; z_correct<="1110111000001000";
        when 7343 => y_in <= "10011100"; x_in <= "00101111"; z_correct<="1110110110100100";
        when 7344 => y_in <= "10011100"; x_in <= "00110000"; z_correct<="1110110101000000";
        when 7345 => y_in <= "10011100"; x_in <= "00110001"; z_correct<="1110110011011100";
        when 7346 => y_in <= "10011100"; x_in <= "00110010"; z_correct<="1110110001111000";
        when 7347 => y_in <= "10011100"; x_in <= "00110011"; z_correct<="1110110000010100";
        when 7348 => y_in <= "10011100"; x_in <= "00110100"; z_correct<="1110101110110000";
        when 7349 => y_in <= "10011100"; x_in <= "00110101"; z_correct<="1110101101001100";
        when 7350 => y_in <= "10011100"; x_in <= "00110110"; z_correct<="1110101011101000";
        when 7351 => y_in <= "10011100"; x_in <= "00110111"; z_correct<="1110101010000100";
        when 7352 => y_in <= "10011100"; x_in <= "00111000"; z_correct<="1110101000100000";
        when 7353 => y_in <= "10011100"; x_in <= "00111001"; z_correct<="1110100110111100";
        when 7354 => y_in <= "10011100"; x_in <= "00111010"; z_correct<="1110100101011000";
        when 7355 => y_in <= "10011100"; x_in <= "00111011"; z_correct<="1110100011110100";
        when 7356 => y_in <= "10011100"; x_in <= "00111100"; z_correct<="1110100010010000";
        when 7357 => y_in <= "10011100"; x_in <= "00111101"; z_correct<="1110100000101100";
        when 7358 => y_in <= "10011100"; x_in <= "00111110"; z_correct<="1110011111001000";
        when 7359 => y_in <= "10011100"; x_in <= "00111111"; z_correct<="1110011101100100";
        when 7360 => y_in <= "10011100"; x_in <= "01000000"; z_correct<="1110011100000000";
        when 7361 => y_in <= "10011100"; x_in <= "01000001"; z_correct<="1110011010011100";
        when 7362 => y_in <= "10011100"; x_in <= "01000010"; z_correct<="1110011000111000";
        when 7363 => y_in <= "10011100"; x_in <= "01000011"; z_correct<="1110010111010100";
        when 7364 => y_in <= "10011100"; x_in <= "01000100"; z_correct<="1110010101110000";
        when 7365 => y_in <= "10011100"; x_in <= "01000101"; z_correct<="1110010100001100";
        when 7366 => y_in <= "10011100"; x_in <= "01000110"; z_correct<="1110010010101000";
        when 7367 => y_in <= "10011100"; x_in <= "01000111"; z_correct<="1110010001000100";
        when 7368 => y_in <= "10011100"; x_in <= "01001000"; z_correct<="1110001111100000";
        when 7369 => y_in <= "10011100"; x_in <= "01001001"; z_correct<="1110001101111100";
        when 7370 => y_in <= "10011100"; x_in <= "01001010"; z_correct<="1110001100011000";
        when 7371 => y_in <= "10011100"; x_in <= "01001011"; z_correct<="1110001010110100";
        when 7372 => y_in <= "10011100"; x_in <= "01001100"; z_correct<="1110001001010000";
        when 7373 => y_in <= "10011100"; x_in <= "01001101"; z_correct<="1110000111101100";
        when 7374 => y_in <= "10011100"; x_in <= "01001110"; z_correct<="1110000110001000";
        when 7375 => y_in <= "10011100"; x_in <= "01001111"; z_correct<="1110000100100100";
        when 7376 => y_in <= "10011100"; x_in <= "01010000"; z_correct<="1110000011000000";
        when 7377 => y_in <= "10011100"; x_in <= "01010001"; z_correct<="1110000001011100";
        when 7378 => y_in <= "10011100"; x_in <= "01010010"; z_correct<="1101111111111000";
        when 7379 => y_in <= "10011100"; x_in <= "01010011"; z_correct<="1101111110010100";
        when 7380 => y_in <= "10011100"; x_in <= "01010100"; z_correct<="1101111100110000";
        when 7381 => y_in <= "10011100"; x_in <= "01010101"; z_correct<="1101111011001100";
        when 7382 => y_in <= "10011100"; x_in <= "01010110"; z_correct<="1101111001101000";
        when 7383 => y_in <= "10011100"; x_in <= "01010111"; z_correct<="1101111000000100";
        when 7384 => y_in <= "10011100"; x_in <= "01011000"; z_correct<="1101110110100000";
        when 7385 => y_in <= "10011100"; x_in <= "01011001"; z_correct<="1101110100111100";
        when 7386 => y_in <= "10011100"; x_in <= "01011010"; z_correct<="1101110011011000";
        when 7387 => y_in <= "10011100"; x_in <= "01011011"; z_correct<="1101110001110100";
        when 7388 => y_in <= "10011100"; x_in <= "01011100"; z_correct<="1101110000010000";
        when 7389 => y_in <= "10011100"; x_in <= "01011101"; z_correct<="1101101110101100";
        when 7390 => y_in <= "10011100"; x_in <= "01011110"; z_correct<="1101101101001000";
        when 7391 => y_in <= "10011100"; x_in <= "01011111"; z_correct<="1101101011100100";
        when 7392 => y_in <= "10011100"; x_in <= "01100000"; z_correct<="1101101010000000";
        when 7393 => y_in <= "10011100"; x_in <= "01100001"; z_correct<="1101101000011100";
        when 7394 => y_in <= "10011100"; x_in <= "01100010"; z_correct<="1101100110111000";
        when 7395 => y_in <= "10011100"; x_in <= "01100011"; z_correct<="1101100101010100";
        when 7396 => y_in <= "10011100"; x_in <= "01100100"; z_correct<="1101100011110000";
        when 7397 => y_in <= "10011100"; x_in <= "01100101"; z_correct<="1101100010001100";
        when 7398 => y_in <= "10011100"; x_in <= "01100110"; z_correct<="1101100000101000";
        when 7399 => y_in <= "10011100"; x_in <= "01100111"; z_correct<="1101011111000100";
        when 7400 => y_in <= "10011100"; x_in <= "01101000"; z_correct<="1101011101100000";
        when 7401 => y_in <= "10011100"; x_in <= "01101001"; z_correct<="1101011011111100";
        when 7402 => y_in <= "10011100"; x_in <= "01101010"; z_correct<="1101011010011000";
        when 7403 => y_in <= "10011100"; x_in <= "01101011"; z_correct<="1101011000110100";
        when 7404 => y_in <= "10011100"; x_in <= "01101100"; z_correct<="1101010111010000";
        when 7405 => y_in <= "10011100"; x_in <= "01101101"; z_correct<="1101010101101100";
        when 7406 => y_in <= "10011100"; x_in <= "01101110"; z_correct<="1101010100001000";
        when 7407 => y_in <= "10011100"; x_in <= "01101111"; z_correct<="1101010010100100";
        when 7408 => y_in <= "10011100"; x_in <= "01110000"; z_correct<="1101010001000000";
        when 7409 => y_in <= "10011100"; x_in <= "01110001"; z_correct<="1101001111011100";
        when 7410 => y_in <= "10011100"; x_in <= "01110010"; z_correct<="1101001101111000";
        when 7411 => y_in <= "10011100"; x_in <= "01110011"; z_correct<="1101001100010100";
        when 7412 => y_in <= "10011100"; x_in <= "01110100"; z_correct<="1101001010110000";
        when 7413 => y_in <= "10011100"; x_in <= "01110101"; z_correct<="1101001001001100";
        when 7414 => y_in <= "10011100"; x_in <= "01110110"; z_correct<="1101000111101000";
        when 7415 => y_in <= "10011100"; x_in <= "01110111"; z_correct<="1101000110000100";
        when 7416 => y_in <= "10011100"; x_in <= "01111000"; z_correct<="1101000100100000";
        when 7417 => y_in <= "10011100"; x_in <= "01111001"; z_correct<="1101000010111100";
        when 7418 => y_in <= "10011100"; x_in <= "01111010"; z_correct<="1101000001011000";
        when 7419 => y_in <= "10011100"; x_in <= "01111011"; z_correct<="1100111111110100";
        when 7420 => y_in <= "10011100"; x_in <= "01111100"; z_correct<="1100111110010000";
        when 7421 => y_in <= "10011100"; x_in <= "01111101"; z_correct<="1100111100101100";
        when 7422 => y_in <= "10011100"; x_in <= "01111110"; z_correct<="1100111011001000";
        when 7423 => y_in <= "10011100"; x_in <= "01111111"; z_correct<="1100111001100100";
        when 7424 => y_in <= "10011101"; x_in <= "10000000"; z_correct<="0011000110000000";
        when 7425 => y_in <= "10011101"; x_in <= "10000001"; z_correct<="0011000100011101";
        when 7426 => y_in <= "10011101"; x_in <= "10000010"; z_correct<="0011000010111010";
        when 7427 => y_in <= "10011101"; x_in <= "10000011"; z_correct<="0011000001010111";
        when 7428 => y_in <= "10011101"; x_in <= "10000100"; z_correct<="0010111111110100";
        when 7429 => y_in <= "10011101"; x_in <= "10000101"; z_correct<="0010111110010001";
        when 7430 => y_in <= "10011101"; x_in <= "10000110"; z_correct<="0010111100101110";
        when 7431 => y_in <= "10011101"; x_in <= "10000111"; z_correct<="0010111011001011";
        when 7432 => y_in <= "10011101"; x_in <= "10001000"; z_correct<="0010111001101000";
        when 7433 => y_in <= "10011101"; x_in <= "10001001"; z_correct<="0010111000000101";
        when 7434 => y_in <= "10011101"; x_in <= "10001010"; z_correct<="0010110110100010";
        when 7435 => y_in <= "10011101"; x_in <= "10001011"; z_correct<="0010110100111111";
        when 7436 => y_in <= "10011101"; x_in <= "10001100"; z_correct<="0010110011011100";
        when 7437 => y_in <= "10011101"; x_in <= "10001101"; z_correct<="0010110001111001";
        when 7438 => y_in <= "10011101"; x_in <= "10001110"; z_correct<="0010110000010110";
        when 7439 => y_in <= "10011101"; x_in <= "10001111"; z_correct<="0010101110110011";
        when 7440 => y_in <= "10011101"; x_in <= "10010000"; z_correct<="0010101101010000";
        when 7441 => y_in <= "10011101"; x_in <= "10010001"; z_correct<="0010101011101101";
        when 7442 => y_in <= "10011101"; x_in <= "10010010"; z_correct<="0010101010001010";
        when 7443 => y_in <= "10011101"; x_in <= "10010011"; z_correct<="0010101000100111";
        when 7444 => y_in <= "10011101"; x_in <= "10010100"; z_correct<="0010100111000100";
        when 7445 => y_in <= "10011101"; x_in <= "10010101"; z_correct<="0010100101100001";
        when 7446 => y_in <= "10011101"; x_in <= "10010110"; z_correct<="0010100011111110";
        when 7447 => y_in <= "10011101"; x_in <= "10010111"; z_correct<="0010100010011011";
        when 7448 => y_in <= "10011101"; x_in <= "10011000"; z_correct<="0010100000111000";
        when 7449 => y_in <= "10011101"; x_in <= "10011001"; z_correct<="0010011111010101";
        when 7450 => y_in <= "10011101"; x_in <= "10011010"; z_correct<="0010011101110010";
        when 7451 => y_in <= "10011101"; x_in <= "10011011"; z_correct<="0010011100001111";
        when 7452 => y_in <= "10011101"; x_in <= "10011100"; z_correct<="0010011010101100";
        when 7453 => y_in <= "10011101"; x_in <= "10011101"; z_correct<="0010011001001001";
        when 7454 => y_in <= "10011101"; x_in <= "10011110"; z_correct<="0010010111100110";
        when 7455 => y_in <= "10011101"; x_in <= "10011111"; z_correct<="0010010110000011";
        when 7456 => y_in <= "10011101"; x_in <= "10100000"; z_correct<="0010010100100000";
        when 7457 => y_in <= "10011101"; x_in <= "10100001"; z_correct<="0010010010111101";
        when 7458 => y_in <= "10011101"; x_in <= "10100010"; z_correct<="0010010001011010";
        when 7459 => y_in <= "10011101"; x_in <= "10100011"; z_correct<="0010001111110111";
        when 7460 => y_in <= "10011101"; x_in <= "10100100"; z_correct<="0010001110010100";
        when 7461 => y_in <= "10011101"; x_in <= "10100101"; z_correct<="0010001100110001";
        when 7462 => y_in <= "10011101"; x_in <= "10100110"; z_correct<="0010001011001110";
        when 7463 => y_in <= "10011101"; x_in <= "10100111"; z_correct<="0010001001101011";
        when 7464 => y_in <= "10011101"; x_in <= "10101000"; z_correct<="0010001000001000";
        when 7465 => y_in <= "10011101"; x_in <= "10101001"; z_correct<="0010000110100101";
        when 7466 => y_in <= "10011101"; x_in <= "10101010"; z_correct<="0010000101000010";
        when 7467 => y_in <= "10011101"; x_in <= "10101011"; z_correct<="0010000011011111";
        when 7468 => y_in <= "10011101"; x_in <= "10101100"; z_correct<="0010000001111100";
        when 7469 => y_in <= "10011101"; x_in <= "10101101"; z_correct<="0010000000011001";
        when 7470 => y_in <= "10011101"; x_in <= "10101110"; z_correct<="0001111110110110";
        when 7471 => y_in <= "10011101"; x_in <= "10101111"; z_correct<="0001111101010011";
        when 7472 => y_in <= "10011101"; x_in <= "10110000"; z_correct<="0001111011110000";
        when 7473 => y_in <= "10011101"; x_in <= "10110001"; z_correct<="0001111010001101";
        when 7474 => y_in <= "10011101"; x_in <= "10110010"; z_correct<="0001111000101010";
        when 7475 => y_in <= "10011101"; x_in <= "10110011"; z_correct<="0001110111000111";
        when 7476 => y_in <= "10011101"; x_in <= "10110100"; z_correct<="0001110101100100";
        when 7477 => y_in <= "10011101"; x_in <= "10110101"; z_correct<="0001110100000001";
        when 7478 => y_in <= "10011101"; x_in <= "10110110"; z_correct<="0001110010011110";
        when 7479 => y_in <= "10011101"; x_in <= "10110111"; z_correct<="0001110000111011";
        when 7480 => y_in <= "10011101"; x_in <= "10111000"; z_correct<="0001101111011000";
        when 7481 => y_in <= "10011101"; x_in <= "10111001"; z_correct<="0001101101110101";
        when 7482 => y_in <= "10011101"; x_in <= "10111010"; z_correct<="0001101100010010";
        when 7483 => y_in <= "10011101"; x_in <= "10111011"; z_correct<="0001101010101111";
        when 7484 => y_in <= "10011101"; x_in <= "10111100"; z_correct<="0001101001001100";
        when 7485 => y_in <= "10011101"; x_in <= "10111101"; z_correct<="0001100111101001";
        when 7486 => y_in <= "10011101"; x_in <= "10111110"; z_correct<="0001100110000110";
        when 7487 => y_in <= "10011101"; x_in <= "10111111"; z_correct<="0001100100100011";
        when 7488 => y_in <= "10011101"; x_in <= "11000000"; z_correct<="0001100011000000";
        when 7489 => y_in <= "10011101"; x_in <= "11000001"; z_correct<="0001100001011101";
        when 7490 => y_in <= "10011101"; x_in <= "11000010"; z_correct<="0001011111111010";
        when 7491 => y_in <= "10011101"; x_in <= "11000011"; z_correct<="0001011110010111";
        when 7492 => y_in <= "10011101"; x_in <= "11000100"; z_correct<="0001011100110100";
        when 7493 => y_in <= "10011101"; x_in <= "11000101"; z_correct<="0001011011010001";
        when 7494 => y_in <= "10011101"; x_in <= "11000110"; z_correct<="0001011001101110";
        when 7495 => y_in <= "10011101"; x_in <= "11000111"; z_correct<="0001011000001011";
        when 7496 => y_in <= "10011101"; x_in <= "11001000"; z_correct<="0001010110101000";
        when 7497 => y_in <= "10011101"; x_in <= "11001001"; z_correct<="0001010101000101";
        when 7498 => y_in <= "10011101"; x_in <= "11001010"; z_correct<="0001010011100010";
        when 7499 => y_in <= "10011101"; x_in <= "11001011"; z_correct<="0001010001111111";
        when 7500 => y_in <= "10011101"; x_in <= "11001100"; z_correct<="0001010000011100";
        when 7501 => y_in <= "10011101"; x_in <= "11001101"; z_correct<="0001001110111001";
        when 7502 => y_in <= "10011101"; x_in <= "11001110"; z_correct<="0001001101010110";
        when 7503 => y_in <= "10011101"; x_in <= "11001111"; z_correct<="0001001011110011";
        when 7504 => y_in <= "10011101"; x_in <= "11010000"; z_correct<="0001001010010000";
        when 7505 => y_in <= "10011101"; x_in <= "11010001"; z_correct<="0001001000101101";
        when 7506 => y_in <= "10011101"; x_in <= "11010010"; z_correct<="0001000111001010";
        when 7507 => y_in <= "10011101"; x_in <= "11010011"; z_correct<="0001000101100111";
        when 7508 => y_in <= "10011101"; x_in <= "11010100"; z_correct<="0001000100000100";
        when 7509 => y_in <= "10011101"; x_in <= "11010101"; z_correct<="0001000010100001";
        when 7510 => y_in <= "10011101"; x_in <= "11010110"; z_correct<="0001000000111110";
        when 7511 => y_in <= "10011101"; x_in <= "11010111"; z_correct<="0000111111011011";
        when 7512 => y_in <= "10011101"; x_in <= "11011000"; z_correct<="0000111101111000";
        when 7513 => y_in <= "10011101"; x_in <= "11011001"; z_correct<="0000111100010101";
        when 7514 => y_in <= "10011101"; x_in <= "11011010"; z_correct<="0000111010110010";
        when 7515 => y_in <= "10011101"; x_in <= "11011011"; z_correct<="0000111001001111";
        when 7516 => y_in <= "10011101"; x_in <= "11011100"; z_correct<="0000110111101100";
        when 7517 => y_in <= "10011101"; x_in <= "11011101"; z_correct<="0000110110001001";
        when 7518 => y_in <= "10011101"; x_in <= "11011110"; z_correct<="0000110100100110";
        when 7519 => y_in <= "10011101"; x_in <= "11011111"; z_correct<="0000110011000011";
        when 7520 => y_in <= "10011101"; x_in <= "11100000"; z_correct<="0000110001100000";
        when 7521 => y_in <= "10011101"; x_in <= "11100001"; z_correct<="0000101111111101";
        when 7522 => y_in <= "10011101"; x_in <= "11100010"; z_correct<="0000101110011010";
        when 7523 => y_in <= "10011101"; x_in <= "11100011"; z_correct<="0000101100110111";
        when 7524 => y_in <= "10011101"; x_in <= "11100100"; z_correct<="0000101011010100";
        when 7525 => y_in <= "10011101"; x_in <= "11100101"; z_correct<="0000101001110001";
        when 7526 => y_in <= "10011101"; x_in <= "11100110"; z_correct<="0000101000001110";
        when 7527 => y_in <= "10011101"; x_in <= "11100111"; z_correct<="0000100110101011";
        when 7528 => y_in <= "10011101"; x_in <= "11101000"; z_correct<="0000100101001000";
        when 7529 => y_in <= "10011101"; x_in <= "11101001"; z_correct<="0000100011100101";
        when 7530 => y_in <= "10011101"; x_in <= "11101010"; z_correct<="0000100010000010";
        when 7531 => y_in <= "10011101"; x_in <= "11101011"; z_correct<="0000100000011111";
        when 7532 => y_in <= "10011101"; x_in <= "11101100"; z_correct<="0000011110111100";
        when 7533 => y_in <= "10011101"; x_in <= "11101101"; z_correct<="0000011101011001";
        when 7534 => y_in <= "10011101"; x_in <= "11101110"; z_correct<="0000011011110110";
        when 7535 => y_in <= "10011101"; x_in <= "11101111"; z_correct<="0000011010010011";
        when 7536 => y_in <= "10011101"; x_in <= "11110000"; z_correct<="0000011000110000";
        when 7537 => y_in <= "10011101"; x_in <= "11110001"; z_correct<="0000010111001101";
        when 7538 => y_in <= "10011101"; x_in <= "11110010"; z_correct<="0000010101101010";
        when 7539 => y_in <= "10011101"; x_in <= "11110011"; z_correct<="0000010100000111";
        when 7540 => y_in <= "10011101"; x_in <= "11110100"; z_correct<="0000010010100100";
        when 7541 => y_in <= "10011101"; x_in <= "11110101"; z_correct<="0000010001000001";
        when 7542 => y_in <= "10011101"; x_in <= "11110110"; z_correct<="0000001111011110";
        when 7543 => y_in <= "10011101"; x_in <= "11110111"; z_correct<="0000001101111011";
        when 7544 => y_in <= "10011101"; x_in <= "11111000"; z_correct<="0000001100011000";
        when 7545 => y_in <= "10011101"; x_in <= "11111001"; z_correct<="0000001010110101";
        when 7546 => y_in <= "10011101"; x_in <= "11111010"; z_correct<="0000001001010010";
        when 7547 => y_in <= "10011101"; x_in <= "11111011"; z_correct<="0000000111101111";
        when 7548 => y_in <= "10011101"; x_in <= "11111100"; z_correct<="0000000110001100";
        when 7549 => y_in <= "10011101"; x_in <= "11111101"; z_correct<="0000000100101001";
        when 7550 => y_in <= "10011101"; x_in <= "11111110"; z_correct<="0000000011000110";
        when 7551 => y_in <= "10011101"; x_in <= "11111111"; z_correct<="0000000001100011";
        when 7552 => y_in <= "10011101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 7553 => y_in <= "10011101"; x_in <= "00000001"; z_correct<="1111111110011101";
        when 7554 => y_in <= "10011101"; x_in <= "00000010"; z_correct<="1111111100111010";
        when 7555 => y_in <= "10011101"; x_in <= "00000011"; z_correct<="1111111011010111";
        when 7556 => y_in <= "10011101"; x_in <= "00000100"; z_correct<="1111111001110100";
        when 7557 => y_in <= "10011101"; x_in <= "00000101"; z_correct<="1111111000010001";
        when 7558 => y_in <= "10011101"; x_in <= "00000110"; z_correct<="1111110110101110";
        when 7559 => y_in <= "10011101"; x_in <= "00000111"; z_correct<="1111110101001011";
        when 7560 => y_in <= "10011101"; x_in <= "00001000"; z_correct<="1111110011101000";
        when 7561 => y_in <= "10011101"; x_in <= "00001001"; z_correct<="1111110010000101";
        when 7562 => y_in <= "10011101"; x_in <= "00001010"; z_correct<="1111110000100010";
        when 7563 => y_in <= "10011101"; x_in <= "00001011"; z_correct<="1111101110111111";
        when 7564 => y_in <= "10011101"; x_in <= "00001100"; z_correct<="1111101101011100";
        when 7565 => y_in <= "10011101"; x_in <= "00001101"; z_correct<="1111101011111001";
        when 7566 => y_in <= "10011101"; x_in <= "00001110"; z_correct<="1111101010010110";
        when 7567 => y_in <= "10011101"; x_in <= "00001111"; z_correct<="1111101000110011";
        when 7568 => y_in <= "10011101"; x_in <= "00010000"; z_correct<="1111100111010000";
        when 7569 => y_in <= "10011101"; x_in <= "00010001"; z_correct<="1111100101101101";
        when 7570 => y_in <= "10011101"; x_in <= "00010010"; z_correct<="1111100100001010";
        when 7571 => y_in <= "10011101"; x_in <= "00010011"; z_correct<="1111100010100111";
        when 7572 => y_in <= "10011101"; x_in <= "00010100"; z_correct<="1111100001000100";
        when 7573 => y_in <= "10011101"; x_in <= "00010101"; z_correct<="1111011111100001";
        when 7574 => y_in <= "10011101"; x_in <= "00010110"; z_correct<="1111011101111110";
        when 7575 => y_in <= "10011101"; x_in <= "00010111"; z_correct<="1111011100011011";
        when 7576 => y_in <= "10011101"; x_in <= "00011000"; z_correct<="1111011010111000";
        when 7577 => y_in <= "10011101"; x_in <= "00011001"; z_correct<="1111011001010101";
        when 7578 => y_in <= "10011101"; x_in <= "00011010"; z_correct<="1111010111110010";
        when 7579 => y_in <= "10011101"; x_in <= "00011011"; z_correct<="1111010110001111";
        when 7580 => y_in <= "10011101"; x_in <= "00011100"; z_correct<="1111010100101100";
        when 7581 => y_in <= "10011101"; x_in <= "00011101"; z_correct<="1111010011001001";
        when 7582 => y_in <= "10011101"; x_in <= "00011110"; z_correct<="1111010001100110";
        when 7583 => y_in <= "10011101"; x_in <= "00011111"; z_correct<="1111010000000011";
        when 7584 => y_in <= "10011101"; x_in <= "00100000"; z_correct<="1111001110100000";
        when 7585 => y_in <= "10011101"; x_in <= "00100001"; z_correct<="1111001100111101";
        when 7586 => y_in <= "10011101"; x_in <= "00100010"; z_correct<="1111001011011010";
        when 7587 => y_in <= "10011101"; x_in <= "00100011"; z_correct<="1111001001110111";
        when 7588 => y_in <= "10011101"; x_in <= "00100100"; z_correct<="1111001000010100";
        when 7589 => y_in <= "10011101"; x_in <= "00100101"; z_correct<="1111000110110001";
        when 7590 => y_in <= "10011101"; x_in <= "00100110"; z_correct<="1111000101001110";
        when 7591 => y_in <= "10011101"; x_in <= "00100111"; z_correct<="1111000011101011";
        when 7592 => y_in <= "10011101"; x_in <= "00101000"; z_correct<="1111000010001000";
        when 7593 => y_in <= "10011101"; x_in <= "00101001"; z_correct<="1111000000100101";
        when 7594 => y_in <= "10011101"; x_in <= "00101010"; z_correct<="1110111111000010";
        when 7595 => y_in <= "10011101"; x_in <= "00101011"; z_correct<="1110111101011111";
        when 7596 => y_in <= "10011101"; x_in <= "00101100"; z_correct<="1110111011111100";
        when 7597 => y_in <= "10011101"; x_in <= "00101101"; z_correct<="1110111010011001";
        when 7598 => y_in <= "10011101"; x_in <= "00101110"; z_correct<="1110111000110110";
        when 7599 => y_in <= "10011101"; x_in <= "00101111"; z_correct<="1110110111010011";
        when 7600 => y_in <= "10011101"; x_in <= "00110000"; z_correct<="1110110101110000";
        when 7601 => y_in <= "10011101"; x_in <= "00110001"; z_correct<="1110110100001101";
        when 7602 => y_in <= "10011101"; x_in <= "00110010"; z_correct<="1110110010101010";
        when 7603 => y_in <= "10011101"; x_in <= "00110011"; z_correct<="1110110001000111";
        when 7604 => y_in <= "10011101"; x_in <= "00110100"; z_correct<="1110101111100100";
        when 7605 => y_in <= "10011101"; x_in <= "00110101"; z_correct<="1110101110000001";
        when 7606 => y_in <= "10011101"; x_in <= "00110110"; z_correct<="1110101100011110";
        when 7607 => y_in <= "10011101"; x_in <= "00110111"; z_correct<="1110101010111011";
        when 7608 => y_in <= "10011101"; x_in <= "00111000"; z_correct<="1110101001011000";
        when 7609 => y_in <= "10011101"; x_in <= "00111001"; z_correct<="1110100111110101";
        when 7610 => y_in <= "10011101"; x_in <= "00111010"; z_correct<="1110100110010010";
        when 7611 => y_in <= "10011101"; x_in <= "00111011"; z_correct<="1110100100101111";
        when 7612 => y_in <= "10011101"; x_in <= "00111100"; z_correct<="1110100011001100";
        when 7613 => y_in <= "10011101"; x_in <= "00111101"; z_correct<="1110100001101001";
        when 7614 => y_in <= "10011101"; x_in <= "00111110"; z_correct<="1110100000000110";
        when 7615 => y_in <= "10011101"; x_in <= "00111111"; z_correct<="1110011110100011";
        when 7616 => y_in <= "10011101"; x_in <= "01000000"; z_correct<="1110011101000000";
        when 7617 => y_in <= "10011101"; x_in <= "01000001"; z_correct<="1110011011011101";
        when 7618 => y_in <= "10011101"; x_in <= "01000010"; z_correct<="1110011001111010";
        when 7619 => y_in <= "10011101"; x_in <= "01000011"; z_correct<="1110011000010111";
        when 7620 => y_in <= "10011101"; x_in <= "01000100"; z_correct<="1110010110110100";
        when 7621 => y_in <= "10011101"; x_in <= "01000101"; z_correct<="1110010101010001";
        when 7622 => y_in <= "10011101"; x_in <= "01000110"; z_correct<="1110010011101110";
        when 7623 => y_in <= "10011101"; x_in <= "01000111"; z_correct<="1110010010001011";
        when 7624 => y_in <= "10011101"; x_in <= "01001000"; z_correct<="1110010000101000";
        when 7625 => y_in <= "10011101"; x_in <= "01001001"; z_correct<="1110001111000101";
        when 7626 => y_in <= "10011101"; x_in <= "01001010"; z_correct<="1110001101100010";
        when 7627 => y_in <= "10011101"; x_in <= "01001011"; z_correct<="1110001011111111";
        when 7628 => y_in <= "10011101"; x_in <= "01001100"; z_correct<="1110001010011100";
        when 7629 => y_in <= "10011101"; x_in <= "01001101"; z_correct<="1110001000111001";
        when 7630 => y_in <= "10011101"; x_in <= "01001110"; z_correct<="1110000111010110";
        when 7631 => y_in <= "10011101"; x_in <= "01001111"; z_correct<="1110000101110011";
        when 7632 => y_in <= "10011101"; x_in <= "01010000"; z_correct<="1110000100010000";
        when 7633 => y_in <= "10011101"; x_in <= "01010001"; z_correct<="1110000010101101";
        when 7634 => y_in <= "10011101"; x_in <= "01010010"; z_correct<="1110000001001010";
        when 7635 => y_in <= "10011101"; x_in <= "01010011"; z_correct<="1101111111100111";
        when 7636 => y_in <= "10011101"; x_in <= "01010100"; z_correct<="1101111110000100";
        when 7637 => y_in <= "10011101"; x_in <= "01010101"; z_correct<="1101111100100001";
        when 7638 => y_in <= "10011101"; x_in <= "01010110"; z_correct<="1101111010111110";
        when 7639 => y_in <= "10011101"; x_in <= "01010111"; z_correct<="1101111001011011";
        when 7640 => y_in <= "10011101"; x_in <= "01011000"; z_correct<="1101110111111000";
        when 7641 => y_in <= "10011101"; x_in <= "01011001"; z_correct<="1101110110010101";
        when 7642 => y_in <= "10011101"; x_in <= "01011010"; z_correct<="1101110100110010";
        when 7643 => y_in <= "10011101"; x_in <= "01011011"; z_correct<="1101110011001111";
        when 7644 => y_in <= "10011101"; x_in <= "01011100"; z_correct<="1101110001101100";
        when 7645 => y_in <= "10011101"; x_in <= "01011101"; z_correct<="1101110000001001";
        when 7646 => y_in <= "10011101"; x_in <= "01011110"; z_correct<="1101101110100110";
        when 7647 => y_in <= "10011101"; x_in <= "01011111"; z_correct<="1101101101000011";
        when 7648 => y_in <= "10011101"; x_in <= "01100000"; z_correct<="1101101011100000";
        when 7649 => y_in <= "10011101"; x_in <= "01100001"; z_correct<="1101101001111101";
        when 7650 => y_in <= "10011101"; x_in <= "01100010"; z_correct<="1101101000011010";
        when 7651 => y_in <= "10011101"; x_in <= "01100011"; z_correct<="1101100110110111";
        when 7652 => y_in <= "10011101"; x_in <= "01100100"; z_correct<="1101100101010100";
        when 7653 => y_in <= "10011101"; x_in <= "01100101"; z_correct<="1101100011110001";
        when 7654 => y_in <= "10011101"; x_in <= "01100110"; z_correct<="1101100010001110";
        when 7655 => y_in <= "10011101"; x_in <= "01100111"; z_correct<="1101100000101011";
        when 7656 => y_in <= "10011101"; x_in <= "01101000"; z_correct<="1101011111001000";
        when 7657 => y_in <= "10011101"; x_in <= "01101001"; z_correct<="1101011101100101";
        when 7658 => y_in <= "10011101"; x_in <= "01101010"; z_correct<="1101011100000010";
        when 7659 => y_in <= "10011101"; x_in <= "01101011"; z_correct<="1101011010011111";
        when 7660 => y_in <= "10011101"; x_in <= "01101100"; z_correct<="1101011000111100";
        when 7661 => y_in <= "10011101"; x_in <= "01101101"; z_correct<="1101010111011001";
        when 7662 => y_in <= "10011101"; x_in <= "01101110"; z_correct<="1101010101110110";
        when 7663 => y_in <= "10011101"; x_in <= "01101111"; z_correct<="1101010100010011";
        when 7664 => y_in <= "10011101"; x_in <= "01110000"; z_correct<="1101010010110000";
        when 7665 => y_in <= "10011101"; x_in <= "01110001"; z_correct<="1101010001001101";
        when 7666 => y_in <= "10011101"; x_in <= "01110010"; z_correct<="1101001111101010";
        when 7667 => y_in <= "10011101"; x_in <= "01110011"; z_correct<="1101001110000111";
        when 7668 => y_in <= "10011101"; x_in <= "01110100"; z_correct<="1101001100100100";
        when 7669 => y_in <= "10011101"; x_in <= "01110101"; z_correct<="1101001011000001";
        when 7670 => y_in <= "10011101"; x_in <= "01110110"; z_correct<="1101001001011110";
        when 7671 => y_in <= "10011101"; x_in <= "01110111"; z_correct<="1101000111111011";
        when 7672 => y_in <= "10011101"; x_in <= "01111000"; z_correct<="1101000110011000";
        when 7673 => y_in <= "10011101"; x_in <= "01111001"; z_correct<="1101000100110101";
        when 7674 => y_in <= "10011101"; x_in <= "01111010"; z_correct<="1101000011010010";
        when 7675 => y_in <= "10011101"; x_in <= "01111011"; z_correct<="1101000001101111";
        when 7676 => y_in <= "10011101"; x_in <= "01111100"; z_correct<="1101000000001100";
        when 7677 => y_in <= "10011101"; x_in <= "01111101"; z_correct<="1100111110101001";
        when 7678 => y_in <= "10011101"; x_in <= "01111110"; z_correct<="1100111101000110";
        when 7679 => y_in <= "10011101"; x_in <= "01111111"; z_correct<="1100111011100011";
        when 7680 => y_in <= "10011110"; x_in <= "10000000"; z_correct<="0011000100000000";
        when 7681 => y_in <= "10011110"; x_in <= "10000001"; z_correct<="0011000010011110";
        when 7682 => y_in <= "10011110"; x_in <= "10000010"; z_correct<="0011000000111100";
        when 7683 => y_in <= "10011110"; x_in <= "10000011"; z_correct<="0010111111011010";
        when 7684 => y_in <= "10011110"; x_in <= "10000100"; z_correct<="0010111101111000";
        when 7685 => y_in <= "10011110"; x_in <= "10000101"; z_correct<="0010111100010110";
        when 7686 => y_in <= "10011110"; x_in <= "10000110"; z_correct<="0010111010110100";
        when 7687 => y_in <= "10011110"; x_in <= "10000111"; z_correct<="0010111001010010";
        when 7688 => y_in <= "10011110"; x_in <= "10001000"; z_correct<="0010110111110000";
        when 7689 => y_in <= "10011110"; x_in <= "10001001"; z_correct<="0010110110001110";
        when 7690 => y_in <= "10011110"; x_in <= "10001010"; z_correct<="0010110100101100";
        when 7691 => y_in <= "10011110"; x_in <= "10001011"; z_correct<="0010110011001010";
        when 7692 => y_in <= "10011110"; x_in <= "10001100"; z_correct<="0010110001101000";
        when 7693 => y_in <= "10011110"; x_in <= "10001101"; z_correct<="0010110000000110";
        when 7694 => y_in <= "10011110"; x_in <= "10001110"; z_correct<="0010101110100100";
        when 7695 => y_in <= "10011110"; x_in <= "10001111"; z_correct<="0010101101000010";
        when 7696 => y_in <= "10011110"; x_in <= "10010000"; z_correct<="0010101011100000";
        when 7697 => y_in <= "10011110"; x_in <= "10010001"; z_correct<="0010101001111110";
        when 7698 => y_in <= "10011110"; x_in <= "10010010"; z_correct<="0010101000011100";
        when 7699 => y_in <= "10011110"; x_in <= "10010011"; z_correct<="0010100110111010";
        when 7700 => y_in <= "10011110"; x_in <= "10010100"; z_correct<="0010100101011000";
        when 7701 => y_in <= "10011110"; x_in <= "10010101"; z_correct<="0010100011110110";
        when 7702 => y_in <= "10011110"; x_in <= "10010110"; z_correct<="0010100010010100";
        when 7703 => y_in <= "10011110"; x_in <= "10010111"; z_correct<="0010100000110010";
        when 7704 => y_in <= "10011110"; x_in <= "10011000"; z_correct<="0010011111010000";
        when 7705 => y_in <= "10011110"; x_in <= "10011001"; z_correct<="0010011101101110";
        when 7706 => y_in <= "10011110"; x_in <= "10011010"; z_correct<="0010011100001100";
        when 7707 => y_in <= "10011110"; x_in <= "10011011"; z_correct<="0010011010101010";
        when 7708 => y_in <= "10011110"; x_in <= "10011100"; z_correct<="0010011001001000";
        when 7709 => y_in <= "10011110"; x_in <= "10011101"; z_correct<="0010010111100110";
        when 7710 => y_in <= "10011110"; x_in <= "10011110"; z_correct<="0010010110000100";
        when 7711 => y_in <= "10011110"; x_in <= "10011111"; z_correct<="0010010100100010";
        when 7712 => y_in <= "10011110"; x_in <= "10100000"; z_correct<="0010010011000000";
        when 7713 => y_in <= "10011110"; x_in <= "10100001"; z_correct<="0010010001011110";
        when 7714 => y_in <= "10011110"; x_in <= "10100010"; z_correct<="0010001111111100";
        when 7715 => y_in <= "10011110"; x_in <= "10100011"; z_correct<="0010001110011010";
        when 7716 => y_in <= "10011110"; x_in <= "10100100"; z_correct<="0010001100111000";
        when 7717 => y_in <= "10011110"; x_in <= "10100101"; z_correct<="0010001011010110";
        when 7718 => y_in <= "10011110"; x_in <= "10100110"; z_correct<="0010001001110100";
        when 7719 => y_in <= "10011110"; x_in <= "10100111"; z_correct<="0010001000010010";
        when 7720 => y_in <= "10011110"; x_in <= "10101000"; z_correct<="0010000110110000";
        when 7721 => y_in <= "10011110"; x_in <= "10101001"; z_correct<="0010000101001110";
        when 7722 => y_in <= "10011110"; x_in <= "10101010"; z_correct<="0010000011101100";
        when 7723 => y_in <= "10011110"; x_in <= "10101011"; z_correct<="0010000010001010";
        when 7724 => y_in <= "10011110"; x_in <= "10101100"; z_correct<="0010000000101000";
        when 7725 => y_in <= "10011110"; x_in <= "10101101"; z_correct<="0001111111000110";
        when 7726 => y_in <= "10011110"; x_in <= "10101110"; z_correct<="0001111101100100";
        when 7727 => y_in <= "10011110"; x_in <= "10101111"; z_correct<="0001111100000010";
        when 7728 => y_in <= "10011110"; x_in <= "10110000"; z_correct<="0001111010100000";
        when 7729 => y_in <= "10011110"; x_in <= "10110001"; z_correct<="0001111000111110";
        when 7730 => y_in <= "10011110"; x_in <= "10110010"; z_correct<="0001110111011100";
        when 7731 => y_in <= "10011110"; x_in <= "10110011"; z_correct<="0001110101111010";
        when 7732 => y_in <= "10011110"; x_in <= "10110100"; z_correct<="0001110100011000";
        when 7733 => y_in <= "10011110"; x_in <= "10110101"; z_correct<="0001110010110110";
        when 7734 => y_in <= "10011110"; x_in <= "10110110"; z_correct<="0001110001010100";
        when 7735 => y_in <= "10011110"; x_in <= "10110111"; z_correct<="0001101111110010";
        when 7736 => y_in <= "10011110"; x_in <= "10111000"; z_correct<="0001101110010000";
        when 7737 => y_in <= "10011110"; x_in <= "10111001"; z_correct<="0001101100101110";
        when 7738 => y_in <= "10011110"; x_in <= "10111010"; z_correct<="0001101011001100";
        when 7739 => y_in <= "10011110"; x_in <= "10111011"; z_correct<="0001101001101010";
        when 7740 => y_in <= "10011110"; x_in <= "10111100"; z_correct<="0001101000001000";
        when 7741 => y_in <= "10011110"; x_in <= "10111101"; z_correct<="0001100110100110";
        when 7742 => y_in <= "10011110"; x_in <= "10111110"; z_correct<="0001100101000100";
        when 7743 => y_in <= "10011110"; x_in <= "10111111"; z_correct<="0001100011100010";
        when 7744 => y_in <= "10011110"; x_in <= "11000000"; z_correct<="0001100010000000";
        when 7745 => y_in <= "10011110"; x_in <= "11000001"; z_correct<="0001100000011110";
        when 7746 => y_in <= "10011110"; x_in <= "11000010"; z_correct<="0001011110111100";
        when 7747 => y_in <= "10011110"; x_in <= "11000011"; z_correct<="0001011101011010";
        when 7748 => y_in <= "10011110"; x_in <= "11000100"; z_correct<="0001011011111000";
        when 7749 => y_in <= "10011110"; x_in <= "11000101"; z_correct<="0001011010010110";
        when 7750 => y_in <= "10011110"; x_in <= "11000110"; z_correct<="0001011000110100";
        when 7751 => y_in <= "10011110"; x_in <= "11000111"; z_correct<="0001010111010010";
        when 7752 => y_in <= "10011110"; x_in <= "11001000"; z_correct<="0001010101110000";
        when 7753 => y_in <= "10011110"; x_in <= "11001001"; z_correct<="0001010100001110";
        when 7754 => y_in <= "10011110"; x_in <= "11001010"; z_correct<="0001010010101100";
        when 7755 => y_in <= "10011110"; x_in <= "11001011"; z_correct<="0001010001001010";
        when 7756 => y_in <= "10011110"; x_in <= "11001100"; z_correct<="0001001111101000";
        when 7757 => y_in <= "10011110"; x_in <= "11001101"; z_correct<="0001001110000110";
        when 7758 => y_in <= "10011110"; x_in <= "11001110"; z_correct<="0001001100100100";
        when 7759 => y_in <= "10011110"; x_in <= "11001111"; z_correct<="0001001011000010";
        when 7760 => y_in <= "10011110"; x_in <= "11010000"; z_correct<="0001001001100000";
        when 7761 => y_in <= "10011110"; x_in <= "11010001"; z_correct<="0001000111111110";
        when 7762 => y_in <= "10011110"; x_in <= "11010010"; z_correct<="0001000110011100";
        when 7763 => y_in <= "10011110"; x_in <= "11010011"; z_correct<="0001000100111010";
        when 7764 => y_in <= "10011110"; x_in <= "11010100"; z_correct<="0001000011011000";
        when 7765 => y_in <= "10011110"; x_in <= "11010101"; z_correct<="0001000001110110";
        when 7766 => y_in <= "10011110"; x_in <= "11010110"; z_correct<="0001000000010100";
        when 7767 => y_in <= "10011110"; x_in <= "11010111"; z_correct<="0000111110110010";
        when 7768 => y_in <= "10011110"; x_in <= "11011000"; z_correct<="0000111101010000";
        when 7769 => y_in <= "10011110"; x_in <= "11011001"; z_correct<="0000111011101110";
        when 7770 => y_in <= "10011110"; x_in <= "11011010"; z_correct<="0000111010001100";
        when 7771 => y_in <= "10011110"; x_in <= "11011011"; z_correct<="0000111000101010";
        when 7772 => y_in <= "10011110"; x_in <= "11011100"; z_correct<="0000110111001000";
        when 7773 => y_in <= "10011110"; x_in <= "11011101"; z_correct<="0000110101100110";
        when 7774 => y_in <= "10011110"; x_in <= "11011110"; z_correct<="0000110100000100";
        when 7775 => y_in <= "10011110"; x_in <= "11011111"; z_correct<="0000110010100010";
        when 7776 => y_in <= "10011110"; x_in <= "11100000"; z_correct<="0000110001000000";
        when 7777 => y_in <= "10011110"; x_in <= "11100001"; z_correct<="0000101111011110";
        when 7778 => y_in <= "10011110"; x_in <= "11100010"; z_correct<="0000101101111100";
        when 7779 => y_in <= "10011110"; x_in <= "11100011"; z_correct<="0000101100011010";
        when 7780 => y_in <= "10011110"; x_in <= "11100100"; z_correct<="0000101010111000";
        when 7781 => y_in <= "10011110"; x_in <= "11100101"; z_correct<="0000101001010110";
        when 7782 => y_in <= "10011110"; x_in <= "11100110"; z_correct<="0000100111110100";
        when 7783 => y_in <= "10011110"; x_in <= "11100111"; z_correct<="0000100110010010";
        when 7784 => y_in <= "10011110"; x_in <= "11101000"; z_correct<="0000100100110000";
        when 7785 => y_in <= "10011110"; x_in <= "11101001"; z_correct<="0000100011001110";
        when 7786 => y_in <= "10011110"; x_in <= "11101010"; z_correct<="0000100001101100";
        when 7787 => y_in <= "10011110"; x_in <= "11101011"; z_correct<="0000100000001010";
        when 7788 => y_in <= "10011110"; x_in <= "11101100"; z_correct<="0000011110101000";
        when 7789 => y_in <= "10011110"; x_in <= "11101101"; z_correct<="0000011101000110";
        when 7790 => y_in <= "10011110"; x_in <= "11101110"; z_correct<="0000011011100100";
        when 7791 => y_in <= "10011110"; x_in <= "11101111"; z_correct<="0000011010000010";
        when 7792 => y_in <= "10011110"; x_in <= "11110000"; z_correct<="0000011000100000";
        when 7793 => y_in <= "10011110"; x_in <= "11110001"; z_correct<="0000010110111110";
        when 7794 => y_in <= "10011110"; x_in <= "11110010"; z_correct<="0000010101011100";
        when 7795 => y_in <= "10011110"; x_in <= "11110011"; z_correct<="0000010011111010";
        when 7796 => y_in <= "10011110"; x_in <= "11110100"; z_correct<="0000010010011000";
        when 7797 => y_in <= "10011110"; x_in <= "11110101"; z_correct<="0000010000110110";
        when 7798 => y_in <= "10011110"; x_in <= "11110110"; z_correct<="0000001111010100";
        when 7799 => y_in <= "10011110"; x_in <= "11110111"; z_correct<="0000001101110010";
        when 7800 => y_in <= "10011110"; x_in <= "11111000"; z_correct<="0000001100010000";
        when 7801 => y_in <= "10011110"; x_in <= "11111001"; z_correct<="0000001010101110";
        when 7802 => y_in <= "10011110"; x_in <= "11111010"; z_correct<="0000001001001100";
        when 7803 => y_in <= "10011110"; x_in <= "11111011"; z_correct<="0000000111101010";
        when 7804 => y_in <= "10011110"; x_in <= "11111100"; z_correct<="0000000110001000";
        when 7805 => y_in <= "10011110"; x_in <= "11111101"; z_correct<="0000000100100110";
        when 7806 => y_in <= "10011110"; x_in <= "11111110"; z_correct<="0000000011000100";
        when 7807 => y_in <= "10011110"; x_in <= "11111111"; z_correct<="0000000001100010";
        when 7808 => y_in <= "10011110"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 7809 => y_in <= "10011110"; x_in <= "00000001"; z_correct<="1111111110011110";
        when 7810 => y_in <= "10011110"; x_in <= "00000010"; z_correct<="1111111100111100";
        when 7811 => y_in <= "10011110"; x_in <= "00000011"; z_correct<="1111111011011010";
        when 7812 => y_in <= "10011110"; x_in <= "00000100"; z_correct<="1111111001111000";
        when 7813 => y_in <= "10011110"; x_in <= "00000101"; z_correct<="1111111000010110";
        when 7814 => y_in <= "10011110"; x_in <= "00000110"; z_correct<="1111110110110100";
        when 7815 => y_in <= "10011110"; x_in <= "00000111"; z_correct<="1111110101010010";
        when 7816 => y_in <= "10011110"; x_in <= "00001000"; z_correct<="1111110011110000";
        when 7817 => y_in <= "10011110"; x_in <= "00001001"; z_correct<="1111110010001110";
        when 7818 => y_in <= "10011110"; x_in <= "00001010"; z_correct<="1111110000101100";
        when 7819 => y_in <= "10011110"; x_in <= "00001011"; z_correct<="1111101111001010";
        when 7820 => y_in <= "10011110"; x_in <= "00001100"; z_correct<="1111101101101000";
        when 7821 => y_in <= "10011110"; x_in <= "00001101"; z_correct<="1111101100000110";
        when 7822 => y_in <= "10011110"; x_in <= "00001110"; z_correct<="1111101010100100";
        when 7823 => y_in <= "10011110"; x_in <= "00001111"; z_correct<="1111101001000010";
        when 7824 => y_in <= "10011110"; x_in <= "00010000"; z_correct<="1111100111100000";
        when 7825 => y_in <= "10011110"; x_in <= "00010001"; z_correct<="1111100101111110";
        when 7826 => y_in <= "10011110"; x_in <= "00010010"; z_correct<="1111100100011100";
        when 7827 => y_in <= "10011110"; x_in <= "00010011"; z_correct<="1111100010111010";
        when 7828 => y_in <= "10011110"; x_in <= "00010100"; z_correct<="1111100001011000";
        when 7829 => y_in <= "10011110"; x_in <= "00010101"; z_correct<="1111011111110110";
        when 7830 => y_in <= "10011110"; x_in <= "00010110"; z_correct<="1111011110010100";
        when 7831 => y_in <= "10011110"; x_in <= "00010111"; z_correct<="1111011100110010";
        when 7832 => y_in <= "10011110"; x_in <= "00011000"; z_correct<="1111011011010000";
        when 7833 => y_in <= "10011110"; x_in <= "00011001"; z_correct<="1111011001101110";
        when 7834 => y_in <= "10011110"; x_in <= "00011010"; z_correct<="1111011000001100";
        when 7835 => y_in <= "10011110"; x_in <= "00011011"; z_correct<="1111010110101010";
        when 7836 => y_in <= "10011110"; x_in <= "00011100"; z_correct<="1111010101001000";
        when 7837 => y_in <= "10011110"; x_in <= "00011101"; z_correct<="1111010011100110";
        when 7838 => y_in <= "10011110"; x_in <= "00011110"; z_correct<="1111010010000100";
        when 7839 => y_in <= "10011110"; x_in <= "00011111"; z_correct<="1111010000100010";
        when 7840 => y_in <= "10011110"; x_in <= "00100000"; z_correct<="1111001111000000";
        when 7841 => y_in <= "10011110"; x_in <= "00100001"; z_correct<="1111001101011110";
        when 7842 => y_in <= "10011110"; x_in <= "00100010"; z_correct<="1111001011111100";
        when 7843 => y_in <= "10011110"; x_in <= "00100011"; z_correct<="1111001010011010";
        when 7844 => y_in <= "10011110"; x_in <= "00100100"; z_correct<="1111001000111000";
        when 7845 => y_in <= "10011110"; x_in <= "00100101"; z_correct<="1111000111010110";
        when 7846 => y_in <= "10011110"; x_in <= "00100110"; z_correct<="1111000101110100";
        when 7847 => y_in <= "10011110"; x_in <= "00100111"; z_correct<="1111000100010010";
        when 7848 => y_in <= "10011110"; x_in <= "00101000"; z_correct<="1111000010110000";
        when 7849 => y_in <= "10011110"; x_in <= "00101001"; z_correct<="1111000001001110";
        when 7850 => y_in <= "10011110"; x_in <= "00101010"; z_correct<="1110111111101100";
        when 7851 => y_in <= "10011110"; x_in <= "00101011"; z_correct<="1110111110001010";
        when 7852 => y_in <= "10011110"; x_in <= "00101100"; z_correct<="1110111100101000";
        when 7853 => y_in <= "10011110"; x_in <= "00101101"; z_correct<="1110111011000110";
        when 7854 => y_in <= "10011110"; x_in <= "00101110"; z_correct<="1110111001100100";
        when 7855 => y_in <= "10011110"; x_in <= "00101111"; z_correct<="1110111000000010";
        when 7856 => y_in <= "10011110"; x_in <= "00110000"; z_correct<="1110110110100000";
        when 7857 => y_in <= "10011110"; x_in <= "00110001"; z_correct<="1110110100111110";
        when 7858 => y_in <= "10011110"; x_in <= "00110010"; z_correct<="1110110011011100";
        when 7859 => y_in <= "10011110"; x_in <= "00110011"; z_correct<="1110110001111010";
        when 7860 => y_in <= "10011110"; x_in <= "00110100"; z_correct<="1110110000011000";
        when 7861 => y_in <= "10011110"; x_in <= "00110101"; z_correct<="1110101110110110";
        when 7862 => y_in <= "10011110"; x_in <= "00110110"; z_correct<="1110101101010100";
        when 7863 => y_in <= "10011110"; x_in <= "00110111"; z_correct<="1110101011110010";
        when 7864 => y_in <= "10011110"; x_in <= "00111000"; z_correct<="1110101010010000";
        when 7865 => y_in <= "10011110"; x_in <= "00111001"; z_correct<="1110101000101110";
        when 7866 => y_in <= "10011110"; x_in <= "00111010"; z_correct<="1110100111001100";
        when 7867 => y_in <= "10011110"; x_in <= "00111011"; z_correct<="1110100101101010";
        when 7868 => y_in <= "10011110"; x_in <= "00111100"; z_correct<="1110100100001000";
        when 7869 => y_in <= "10011110"; x_in <= "00111101"; z_correct<="1110100010100110";
        when 7870 => y_in <= "10011110"; x_in <= "00111110"; z_correct<="1110100001000100";
        when 7871 => y_in <= "10011110"; x_in <= "00111111"; z_correct<="1110011111100010";
        when 7872 => y_in <= "10011110"; x_in <= "01000000"; z_correct<="1110011110000000";
        when 7873 => y_in <= "10011110"; x_in <= "01000001"; z_correct<="1110011100011110";
        when 7874 => y_in <= "10011110"; x_in <= "01000010"; z_correct<="1110011010111100";
        when 7875 => y_in <= "10011110"; x_in <= "01000011"; z_correct<="1110011001011010";
        when 7876 => y_in <= "10011110"; x_in <= "01000100"; z_correct<="1110010111111000";
        when 7877 => y_in <= "10011110"; x_in <= "01000101"; z_correct<="1110010110010110";
        when 7878 => y_in <= "10011110"; x_in <= "01000110"; z_correct<="1110010100110100";
        when 7879 => y_in <= "10011110"; x_in <= "01000111"; z_correct<="1110010011010010";
        when 7880 => y_in <= "10011110"; x_in <= "01001000"; z_correct<="1110010001110000";
        when 7881 => y_in <= "10011110"; x_in <= "01001001"; z_correct<="1110010000001110";
        when 7882 => y_in <= "10011110"; x_in <= "01001010"; z_correct<="1110001110101100";
        when 7883 => y_in <= "10011110"; x_in <= "01001011"; z_correct<="1110001101001010";
        when 7884 => y_in <= "10011110"; x_in <= "01001100"; z_correct<="1110001011101000";
        when 7885 => y_in <= "10011110"; x_in <= "01001101"; z_correct<="1110001010000110";
        when 7886 => y_in <= "10011110"; x_in <= "01001110"; z_correct<="1110001000100100";
        when 7887 => y_in <= "10011110"; x_in <= "01001111"; z_correct<="1110000111000010";
        when 7888 => y_in <= "10011110"; x_in <= "01010000"; z_correct<="1110000101100000";
        when 7889 => y_in <= "10011110"; x_in <= "01010001"; z_correct<="1110000011111110";
        when 7890 => y_in <= "10011110"; x_in <= "01010010"; z_correct<="1110000010011100";
        when 7891 => y_in <= "10011110"; x_in <= "01010011"; z_correct<="1110000000111010";
        when 7892 => y_in <= "10011110"; x_in <= "01010100"; z_correct<="1101111111011000";
        when 7893 => y_in <= "10011110"; x_in <= "01010101"; z_correct<="1101111101110110";
        when 7894 => y_in <= "10011110"; x_in <= "01010110"; z_correct<="1101111100010100";
        when 7895 => y_in <= "10011110"; x_in <= "01010111"; z_correct<="1101111010110010";
        when 7896 => y_in <= "10011110"; x_in <= "01011000"; z_correct<="1101111001010000";
        when 7897 => y_in <= "10011110"; x_in <= "01011001"; z_correct<="1101110111101110";
        when 7898 => y_in <= "10011110"; x_in <= "01011010"; z_correct<="1101110110001100";
        when 7899 => y_in <= "10011110"; x_in <= "01011011"; z_correct<="1101110100101010";
        when 7900 => y_in <= "10011110"; x_in <= "01011100"; z_correct<="1101110011001000";
        when 7901 => y_in <= "10011110"; x_in <= "01011101"; z_correct<="1101110001100110";
        when 7902 => y_in <= "10011110"; x_in <= "01011110"; z_correct<="1101110000000100";
        when 7903 => y_in <= "10011110"; x_in <= "01011111"; z_correct<="1101101110100010";
        when 7904 => y_in <= "10011110"; x_in <= "01100000"; z_correct<="1101101101000000";
        when 7905 => y_in <= "10011110"; x_in <= "01100001"; z_correct<="1101101011011110";
        when 7906 => y_in <= "10011110"; x_in <= "01100010"; z_correct<="1101101001111100";
        when 7907 => y_in <= "10011110"; x_in <= "01100011"; z_correct<="1101101000011010";
        when 7908 => y_in <= "10011110"; x_in <= "01100100"; z_correct<="1101100110111000";
        when 7909 => y_in <= "10011110"; x_in <= "01100101"; z_correct<="1101100101010110";
        when 7910 => y_in <= "10011110"; x_in <= "01100110"; z_correct<="1101100011110100";
        when 7911 => y_in <= "10011110"; x_in <= "01100111"; z_correct<="1101100010010010";
        when 7912 => y_in <= "10011110"; x_in <= "01101000"; z_correct<="1101100000110000";
        when 7913 => y_in <= "10011110"; x_in <= "01101001"; z_correct<="1101011111001110";
        when 7914 => y_in <= "10011110"; x_in <= "01101010"; z_correct<="1101011101101100";
        when 7915 => y_in <= "10011110"; x_in <= "01101011"; z_correct<="1101011100001010";
        when 7916 => y_in <= "10011110"; x_in <= "01101100"; z_correct<="1101011010101000";
        when 7917 => y_in <= "10011110"; x_in <= "01101101"; z_correct<="1101011001000110";
        when 7918 => y_in <= "10011110"; x_in <= "01101110"; z_correct<="1101010111100100";
        when 7919 => y_in <= "10011110"; x_in <= "01101111"; z_correct<="1101010110000010";
        when 7920 => y_in <= "10011110"; x_in <= "01110000"; z_correct<="1101010100100000";
        when 7921 => y_in <= "10011110"; x_in <= "01110001"; z_correct<="1101010010111110";
        when 7922 => y_in <= "10011110"; x_in <= "01110010"; z_correct<="1101010001011100";
        when 7923 => y_in <= "10011110"; x_in <= "01110011"; z_correct<="1101001111111010";
        when 7924 => y_in <= "10011110"; x_in <= "01110100"; z_correct<="1101001110011000";
        when 7925 => y_in <= "10011110"; x_in <= "01110101"; z_correct<="1101001100110110";
        when 7926 => y_in <= "10011110"; x_in <= "01110110"; z_correct<="1101001011010100";
        when 7927 => y_in <= "10011110"; x_in <= "01110111"; z_correct<="1101001001110010";
        when 7928 => y_in <= "10011110"; x_in <= "01111000"; z_correct<="1101001000010000";
        when 7929 => y_in <= "10011110"; x_in <= "01111001"; z_correct<="1101000110101110";
        when 7930 => y_in <= "10011110"; x_in <= "01111010"; z_correct<="1101000101001100";
        when 7931 => y_in <= "10011110"; x_in <= "01111011"; z_correct<="1101000011101010";
        when 7932 => y_in <= "10011110"; x_in <= "01111100"; z_correct<="1101000010001000";
        when 7933 => y_in <= "10011110"; x_in <= "01111101"; z_correct<="1101000000100110";
        when 7934 => y_in <= "10011110"; x_in <= "01111110"; z_correct<="1100111111000100";
        when 7935 => y_in <= "10011110"; x_in <= "01111111"; z_correct<="1100111101100010";
        when 7936 => y_in <= "10011111"; x_in <= "10000000"; z_correct<="0011000010000000";
        when 7937 => y_in <= "10011111"; x_in <= "10000001"; z_correct<="0011000000011111";
        when 7938 => y_in <= "10011111"; x_in <= "10000010"; z_correct<="0010111110111110";
        when 7939 => y_in <= "10011111"; x_in <= "10000011"; z_correct<="0010111101011101";
        when 7940 => y_in <= "10011111"; x_in <= "10000100"; z_correct<="0010111011111100";
        when 7941 => y_in <= "10011111"; x_in <= "10000101"; z_correct<="0010111010011011";
        when 7942 => y_in <= "10011111"; x_in <= "10000110"; z_correct<="0010111000111010";
        when 7943 => y_in <= "10011111"; x_in <= "10000111"; z_correct<="0010110111011001";
        when 7944 => y_in <= "10011111"; x_in <= "10001000"; z_correct<="0010110101111000";
        when 7945 => y_in <= "10011111"; x_in <= "10001001"; z_correct<="0010110100010111";
        when 7946 => y_in <= "10011111"; x_in <= "10001010"; z_correct<="0010110010110110";
        when 7947 => y_in <= "10011111"; x_in <= "10001011"; z_correct<="0010110001010101";
        when 7948 => y_in <= "10011111"; x_in <= "10001100"; z_correct<="0010101111110100";
        when 7949 => y_in <= "10011111"; x_in <= "10001101"; z_correct<="0010101110010011";
        when 7950 => y_in <= "10011111"; x_in <= "10001110"; z_correct<="0010101100110010";
        when 7951 => y_in <= "10011111"; x_in <= "10001111"; z_correct<="0010101011010001";
        when 7952 => y_in <= "10011111"; x_in <= "10010000"; z_correct<="0010101001110000";
        when 7953 => y_in <= "10011111"; x_in <= "10010001"; z_correct<="0010101000001111";
        when 7954 => y_in <= "10011111"; x_in <= "10010010"; z_correct<="0010100110101110";
        when 7955 => y_in <= "10011111"; x_in <= "10010011"; z_correct<="0010100101001101";
        when 7956 => y_in <= "10011111"; x_in <= "10010100"; z_correct<="0010100011101100";
        when 7957 => y_in <= "10011111"; x_in <= "10010101"; z_correct<="0010100010001011";
        when 7958 => y_in <= "10011111"; x_in <= "10010110"; z_correct<="0010100000101010";
        when 7959 => y_in <= "10011111"; x_in <= "10010111"; z_correct<="0010011111001001";
        when 7960 => y_in <= "10011111"; x_in <= "10011000"; z_correct<="0010011101101000";
        when 7961 => y_in <= "10011111"; x_in <= "10011001"; z_correct<="0010011100000111";
        when 7962 => y_in <= "10011111"; x_in <= "10011010"; z_correct<="0010011010100110";
        when 7963 => y_in <= "10011111"; x_in <= "10011011"; z_correct<="0010011001000101";
        when 7964 => y_in <= "10011111"; x_in <= "10011100"; z_correct<="0010010111100100";
        when 7965 => y_in <= "10011111"; x_in <= "10011101"; z_correct<="0010010110000011";
        when 7966 => y_in <= "10011111"; x_in <= "10011110"; z_correct<="0010010100100010";
        when 7967 => y_in <= "10011111"; x_in <= "10011111"; z_correct<="0010010011000001";
        when 7968 => y_in <= "10011111"; x_in <= "10100000"; z_correct<="0010010001100000";
        when 7969 => y_in <= "10011111"; x_in <= "10100001"; z_correct<="0010001111111111";
        when 7970 => y_in <= "10011111"; x_in <= "10100010"; z_correct<="0010001110011110";
        when 7971 => y_in <= "10011111"; x_in <= "10100011"; z_correct<="0010001100111101";
        when 7972 => y_in <= "10011111"; x_in <= "10100100"; z_correct<="0010001011011100";
        when 7973 => y_in <= "10011111"; x_in <= "10100101"; z_correct<="0010001001111011";
        when 7974 => y_in <= "10011111"; x_in <= "10100110"; z_correct<="0010001000011010";
        when 7975 => y_in <= "10011111"; x_in <= "10100111"; z_correct<="0010000110111001";
        when 7976 => y_in <= "10011111"; x_in <= "10101000"; z_correct<="0010000101011000";
        when 7977 => y_in <= "10011111"; x_in <= "10101001"; z_correct<="0010000011110111";
        when 7978 => y_in <= "10011111"; x_in <= "10101010"; z_correct<="0010000010010110";
        when 7979 => y_in <= "10011111"; x_in <= "10101011"; z_correct<="0010000000110101";
        when 7980 => y_in <= "10011111"; x_in <= "10101100"; z_correct<="0001111111010100";
        when 7981 => y_in <= "10011111"; x_in <= "10101101"; z_correct<="0001111101110011";
        when 7982 => y_in <= "10011111"; x_in <= "10101110"; z_correct<="0001111100010010";
        when 7983 => y_in <= "10011111"; x_in <= "10101111"; z_correct<="0001111010110001";
        when 7984 => y_in <= "10011111"; x_in <= "10110000"; z_correct<="0001111001010000";
        when 7985 => y_in <= "10011111"; x_in <= "10110001"; z_correct<="0001110111101111";
        when 7986 => y_in <= "10011111"; x_in <= "10110010"; z_correct<="0001110110001110";
        when 7987 => y_in <= "10011111"; x_in <= "10110011"; z_correct<="0001110100101101";
        when 7988 => y_in <= "10011111"; x_in <= "10110100"; z_correct<="0001110011001100";
        when 7989 => y_in <= "10011111"; x_in <= "10110101"; z_correct<="0001110001101011";
        when 7990 => y_in <= "10011111"; x_in <= "10110110"; z_correct<="0001110000001010";
        when 7991 => y_in <= "10011111"; x_in <= "10110111"; z_correct<="0001101110101001";
        when 7992 => y_in <= "10011111"; x_in <= "10111000"; z_correct<="0001101101001000";
        when 7993 => y_in <= "10011111"; x_in <= "10111001"; z_correct<="0001101011100111";
        when 7994 => y_in <= "10011111"; x_in <= "10111010"; z_correct<="0001101010000110";
        when 7995 => y_in <= "10011111"; x_in <= "10111011"; z_correct<="0001101000100101";
        when 7996 => y_in <= "10011111"; x_in <= "10111100"; z_correct<="0001100111000100";
        when 7997 => y_in <= "10011111"; x_in <= "10111101"; z_correct<="0001100101100011";
        when 7998 => y_in <= "10011111"; x_in <= "10111110"; z_correct<="0001100100000010";
        when 7999 => y_in <= "10011111"; x_in <= "10111111"; z_correct<="0001100010100001";
        when 8000 => y_in <= "10011111"; x_in <= "11000000"; z_correct<="0001100001000000";
        when 8001 => y_in <= "10011111"; x_in <= "11000001"; z_correct<="0001011111011111";
        when 8002 => y_in <= "10011111"; x_in <= "11000010"; z_correct<="0001011101111110";
        when 8003 => y_in <= "10011111"; x_in <= "11000011"; z_correct<="0001011100011101";
        when 8004 => y_in <= "10011111"; x_in <= "11000100"; z_correct<="0001011010111100";
        when 8005 => y_in <= "10011111"; x_in <= "11000101"; z_correct<="0001011001011011";
        when 8006 => y_in <= "10011111"; x_in <= "11000110"; z_correct<="0001010111111010";
        when 8007 => y_in <= "10011111"; x_in <= "11000111"; z_correct<="0001010110011001";
        when 8008 => y_in <= "10011111"; x_in <= "11001000"; z_correct<="0001010100111000";
        when 8009 => y_in <= "10011111"; x_in <= "11001001"; z_correct<="0001010011010111";
        when 8010 => y_in <= "10011111"; x_in <= "11001010"; z_correct<="0001010001110110";
        when 8011 => y_in <= "10011111"; x_in <= "11001011"; z_correct<="0001010000010101";
        when 8012 => y_in <= "10011111"; x_in <= "11001100"; z_correct<="0001001110110100";
        when 8013 => y_in <= "10011111"; x_in <= "11001101"; z_correct<="0001001101010011";
        when 8014 => y_in <= "10011111"; x_in <= "11001110"; z_correct<="0001001011110010";
        when 8015 => y_in <= "10011111"; x_in <= "11001111"; z_correct<="0001001010010001";
        when 8016 => y_in <= "10011111"; x_in <= "11010000"; z_correct<="0001001000110000";
        when 8017 => y_in <= "10011111"; x_in <= "11010001"; z_correct<="0001000111001111";
        when 8018 => y_in <= "10011111"; x_in <= "11010010"; z_correct<="0001000101101110";
        when 8019 => y_in <= "10011111"; x_in <= "11010011"; z_correct<="0001000100001101";
        when 8020 => y_in <= "10011111"; x_in <= "11010100"; z_correct<="0001000010101100";
        when 8021 => y_in <= "10011111"; x_in <= "11010101"; z_correct<="0001000001001011";
        when 8022 => y_in <= "10011111"; x_in <= "11010110"; z_correct<="0000111111101010";
        when 8023 => y_in <= "10011111"; x_in <= "11010111"; z_correct<="0000111110001001";
        when 8024 => y_in <= "10011111"; x_in <= "11011000"; z_correct<="0000111100101000";
        when 8025 => y_in <= "10011111"; x_in <= "11011001"; z_correct<="0000111011000111";
        when 8026 => y_in <= "10011111"; x_in <= "11011010"; z_correct<="0000111001100110";
        when 8027 => y_in <= "10011111"; x_in <= "11011011"; z_correct<="0000111000000101";
        when 8028 => y_in <= "10011111"; x_in <= "11011100"; z_correct<="0000110110100100";
        when 8029 => y_in <= "10011111"; x_in <= "11011101"; z_correct<="0000110101000011";
        when 8030 => y_in <= "10011111"; x_in <= "11011110"; z_correct<="0000110011100010";
        when 8031 => y_in <= "10011111"; x_in <= "11011111"; z_correct<="0000110010000001";
        when 8032 => y_in <= "10011111"; x_in <= "11100000"; z_correct<="0000110000100000";
        when 8033 => y_in <= "10011111"; x_in <= "11100001"; z_correct<="0000101110111111";
        when 8034 => y_in <= "10011111"; x_in <= "11100010"; z_correct<="0000101101011110";
        when 8035 => y_in <= "10011111"; x_in <= "11100011"; z_correct<="0000101011111101";
        when 8036 => y_in <= "10011111"; x_in <= "11100100"; z_correct<="0000101010011100";
        when 8037 => y_in <= "10011111"; x_in <= "11100101"; z_correct<="0000101000111011";
        when 8038 => y_in <= "10011111"; x_in <= "11100110"; z_correct<="0000100111011010";
        when 8039 => y_in <= "10011111"; x_in <= "11100111"; z_correct<="0000100101111001";
        when 8040 => y_in <= "10011111"; x_in <= "11101000"; z_correct<="0000100100011000";
        when 8041 => y_in <= "10011111"; x_in <= "11101001"; z_correct<="0000100010110111";
        when 8042 => y_in <= "10011111"; x_in <= "11101010"; z_correct<="0000100001010110";
        when 8043 => y_in <= "10011111"; x_in <= "11101011"; z_correct<="0000011111110101";
        when 8044 => y_in <= "10011111"; x_in <= "11101100"; z_correct<="0000011110010100";
        when 8045 => y_in <= "10011111"; x_in <= "11101101"; z_correct<="0000011100110011";
        when 8046 => y_in <= "10011111"; x_in <= "11101110"; z_correct<="0000011011010010";
        when 8047 => y_in <= "10011111"; x_in <= "11101111"; z_correct<="0000011001110001";
        when 8048 => y_in <= "10011111"; x_in <= "11110000"; z_correct<="0000011000010000";
        when 8049 => y_in <= "10011111"; x_in <= "11110001"; z_correct<="0000010110101111";
        when 8050 => y_in <= "10011111"; x_in <= "11110010"; z_correct<="0000010101001110";
        when 8051 => y_in <= "10011111"; x_in <= "11110011"; z_correct<="0000010011101101";
        when 8052 => y_in <= "10011111"; x_in <= "11110100"; z_correct<="0000010010001100";
        when 8053 => y_in <= "10011111"; x_in <= "11110101"; z_correct<="0000010000101011";
        when 8054 => y_in <= "10011111"; x_in <= "11110110"; z_correct<="0000001111001010";
        when 8055 => y_in <= "10011111"; x_in <= "11110111"; z_correct<="0000001101101001";
        when 8056 => y_in <= "10011111"; x_in <= "11111000"; z_correct<="0000001100001000";
        when 8057 => y_in <= "10011111"; x_in <= "11111001"; z_correct<="0000001010100111";
        when 8058 => y_in <= "10011111"; x_in <= "11111010"; z_correct<="0000001001000110";
        when 8059 => y_in <= "10011111"; x_in <= "11111011"; z_correct<="0000000111100101";
        when 8060 => y_in <= "10011111"; x_in <= "11111100"; z_correct<="0000000110000100";
        when 8061 => y_in <= "10011111"; x_in <= "11111101"; z_correct<="0000000100100011";
        when 8062 => y_in <= "10011111"; x_in <= "11111110"; z_correct<="0000000011000010";
        when 8063 => y_in <= "10011111"; x_in <= "11111111"; z_correct<="0000000001100001";
        when 8064 => y_in <= "10011111"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 8065 => y_in <= "10011111"; x_in <= "00000001"; z_correct<="1111111110011111";
        when 8066 => y_in <= "10011111"; x_in <= "00000010"; z_correct<="1111111100111110";
        when 8067 => y_in <= "10011111"; x_in <= "00000011"; z_correct<="1111111011011101";
        when 8068 => y_in <= "10011111"; x_in <= "00000100"; z_correct<="1111111001111100";
        when 8069 => y_in <= "10011111"; x_in <= "00000101"; z_correct<="1111111000011011";
        when 8070 => y_in <= "10011111"; x_in <= "00000110"; z_correct<="1111110110111010";
        when 8071 => y_in <= "10011111"; x_in <= "00000111"; z_correct<="1111110101011001";
        when 8072 => y_in <= "10011111"; x_in <= "00001000"; z_correct<="1111110011111000";
        when 8073 => y_in <= "10011111"; x_in <= "00001001"; z_correct<="1111110010010111";
        when 8074 => y_in <= "10011111"; x_in <= "00001010"; z_correct<="1111110000110110";
        when 8075 => y_in <= "10011111"; x_in <= "00001011"; z_correct<="1111101111010101";
        when 8076 => y_in <= "10011111"; x_in <= "00001100"; z_correct<="1111101101110100";
        when 8077 => y_in <= "10011111"; x_in <= "00001101"; z_correct<="1111101100010011";
        when 8078 => y_in <= "10011111"; x_in <= "00001110"; z_correct<="1111101010110010";
        when 8079 => y_in <= "10011111"; x_in <= "00001111"; z_correct<="1111101001010001";
        when 8080 => y_in <= "10011111"; x_in <= "00010000"; z_correct<="1111100111110000";
        when 8081 => y_in <= "10011111"; x_in <= "00010001"; z_correct<="1111100110001111";
        when 8082 => y_in <= "10011111"; x_in <= "00010010"; z_correct<="1111100100101110";
        when 8083 => y_in <= "10011111"; x_in <= "00010011"; z_correct<="1111100011001101";
        when 8084 => y_in <= "10011111"; x_in <= "00010100"; z_correct<="1111100001101100";
        when 8085 => y_in <= "10011111"; x_in <= "00010101"; z_correct<="1111100000001011";
        when 8086 => y_in <= "10011111"; x_in <= "00010110"; z_correct<="1111011110101010";
        when 8087 => y_in <= "10011111"; x_in <= "00010111"; z_correct<="1111011101001001";
        when 8088 => y_in <= "10011111"; x_in <= "00011000"; z_correct<="1111011011101000";
        when 8089 => y_in <= "10011111"; x_in <= "00011001"; z_correct<="1111011010000111";
        when 8090 => y_in <= "10011111"; x_in <= "00011010"; z_correct<="1111011000100110";
        when 8091 => y_in <= "10011111"; x_in <= "00011011"; z_correct<="1111010111000101";
        when 8092 => y_in <= "10011111"; x_in <= "00011100"; z_correct<="1111010101100100";
        when 8093 => y_in <= "10011111"; x_in <= "00011101"; z_correct<="1111010100000011";
        when 8094 => y_in <= "10011111"; x_in <= "00011110"; z_correct<="1111010010100010";
        when 8095 => y_in <= "10011111"; x_in <= "00011111"; z_correct<="1111010001000001";
        when 8096 => y_in <= "10011111"; x_in <= "00100000"; z_correct<="1111001111100000";
        when 8097 => y_in <= "10011111"; x_in <= "00100001"; z_correct<="1111001101111111";
        when 8098 => y_in <= "10011111"; x_in <= "00100010"; z_correct<="1111001100011110";
        when 8099 => y_in <= "10011111"; x_in <= "00100011"; z_correct<="1111001010111101";
        when 8100 => y_in <= "10011111"; x_in <= "00100100"; z_correct<="1111001001011100";
        when 8101 => y_in <= "10011111"; x_in <= "00100101"; z_correct<="1111000111111011";
        when 8102 => y_in <= "10011111"; x_in <= "00100110"; z_correct<="1111000110011010";
        when 8103 => y_in <= "10011111"; x_in <= "00100111"; z_correct<="1111000100111001";
        when 8104 => y_in <= "10011111"; x_in <= "00101000"; z_correct<="1111000011011000";
        when 8105 => y_in <= "10011111"; x_in <= "00101001"; z_correct<="1111000001110111";
        when 8106 => y_in <= "10011111"; x_in <= "00101010"; z_correct<="1111000000010110";
        when 8107 => y_in <= "10011111"; x_in <= "00101011"; z_correct<="1110111110110101";
        when 8108 => y_in <= "10011111"; x_in <= "00101100"; z_correct<="1110111101010100";
        when 8109 => y_in <= "10011111"; x_in <= "00101101"; z_correct<="1110111011110011";
        when 8110 => y_in <= "10011111"; x_in <= "00101110"; z_correct<="1110111010010010";
        when 8111 => y_in <= "10011111"; x_in <= "00101111"; z_correct<="1110111000110001";
        when 8112 => y_in <= "10011111"; x_in <= "00110000"; z_correct<="1110110111010000";
        when 8113 => y_in <= "10011111"; x_in <= "00110001"; z_correct<="1110110101101111";
        when 8114 => y_in <= "10011111"; x_in <= "00110010"; z_correct<="1110110100001110";
        when 8115 => y_in <= "10011111"; x_in <= "00110011"; z_correct<="1110110010101101";
        when 8116 => y_in <= "10011111"; x_in <= "00110100"; z_correct<="1110110001001100";
        when 8117 => y_in <= "10011111"; x_in <= "00110101"; z_correct<="1110101111101011";
        when 8118 => y_in <= "10011111"; x_in <= "00110110"; z_correct<="1110101110001010";
        when 8119 => y_in <= "10011111"; x_in <= "00110111"; z_correct<="1110101100101001";
        when 8120 => y_in <= "10011111"; x_in <= "00111000"; z_correct<="1110101011001000";
        when 8121 => y_in <= "10011111"; x_in <= "00111001"; z_correct<="1110101001100111";
        when 8122 => y_in <= "10011111"; x_in <= "00111010"; z_correct<="1110101000000110";
        when 8123 => y_in <= "10011111"; x_in <= "00111011"; z_correct<="1110100110100101";
        when 8124 => y_in <= "10011111"; x_in <= "00111100"; z_correct<="1110100101000100";
        when 8125 => y_in <= "10011111"; x_in <= "00111101"; z_correct<="1110100011100011";
        when 8126 => y_in <= "10011111"; x_in <= "00111110"; z_correct<="1110100010000010";
        when 8127 => y_in <= "10011111"; x_in <= "00111111"; z_correct<="1110100000100001";
        when 8128 => y_in <= "10011111"; x_in <= "01000000"; z_correct<="1110011111000000";
        when 8129 => y_in <= "10011111"; x_in <= "01000001"; z_correct<="1110011101011111";
        when 8130 => y_in <= "10011111"; x_in <= "01000010"; z_correct<="1110011011111110";
        when 8131 => y_in <= "10011111"; x_in <= "01000011"; z_correct<="1110011010011101";
        when 8132 => y_in <= "10011111"; x_in <= "01000100"; z_correct<="1110011000111100";
        when 8133 => y_in <= "10011111"; x_in <= "01000101"; z_correct<="1110010111011011";
        when 8134 => y_in <= "10011111"; x_in <= "01000110"; z_correct<="1110010101111010";
        when 8135 => y_in <= "10011111"; x_in <= "01000111"; z_correct<="1110010100011001";
        when 8136 => y_in <= "10011111"; x_in <= "01001000"; z_correct<="1110010010111000";
        when 8137 => y_in <= "10011111"; x_in <= "01001001"; z_correct<="1110010001010111";
        when 8138 => y_in <= "10011111"; x_in <= "01001010"; z_correct<="1110001111110110";
        when 8139 => y_in <= "10011111"; x_in <= "01001011"; z_correct<="1110001110010101";
        when 8140 => y_in <= "10011111"; x_in <= "01001100"; z_correct<="1110001100110100";
        when 8141 => y_in <= "10011111"; x_in <= "01001101"; z_correct<="1110001011010011";
        when 8142 => y_in <= "10011111"; x_in <= "01001110"; z_correct<="1110001001110010";
        when 8143 => y_in <= "10011111"; x_in <= "01001111"; z_correct<="1110001000010001";
        when 8144 => y_in <= "10011111"; x_in <= "01010000"; z_correct<="1110000110110000";
        when 8145 => y_in <= "10011111"; x_in <= "01010001"; z_correct<="1110000101001111";
        when 8146 => y_in <= "10011111"; x_in <= "01010010"; z_correct<="1110000011101110";
        when 8147 => y_in <= "10011111"; x_in <= "01010011"; z_correct<="1110000010001101";
        when 8148 => y_in <= "10011111"; x_in <= "01010100"; z_correct<="1110000000101100";
        when 8149 => y_in <= "10011111"; x_in <= "01010101"; z_correct<="1101111111001011";
        when 8150 => y_in <= "10011111"; x_in <= "01010110"; z_correct<="1101111101101010";
        when 8151 => y_in <= "10011111"; x_in <= "01010111"; z_correct<="1101111100001001";
        when 8152 => y_in <= "10011111"; x_in <= "01011000"; z_correct<="1101111010101000";
        when 8153 => y_in <= "10011111"; x_in <= "01011001"; z_correct<="1101111001000111";
        when 8154 => y_in <= "10011111"; x_in <= "01011010"; z_correct<="1101110111100110";
        when 8155 => y_in <= "10011111"; x_in <= "01011011"; z_correct<="1101110110000101";
        when 8156 => y_in <= "10011111"; x_in <= "01011100"; z_correct<="1101110100100100";
        when 8157 => y_in <= "10011111"; x_in <= "01011101"; z_correct<="1101110011000011";
        when 8158 => y_in <= "10011111"; x_in <= "01011110"; z_correct<="1101110001100010";
        when 8159 => y_in <= "10011111"; x_in <= "01011111"; z_correct<="1101110000000001";
        when 8160 => y_in <= "10011111"; x_in <= "01100000"; z_correct<="1101101110100000";
        when 8161 => y_in <= "10011111"; x_in <= "01100001"; z_correct<="1101101100111111";
        when 8162 => y_in <= "10011111"; x_in <= "01100010"; z_correct<="1101101011011110";
        when 8163 => y_in <= "10011111"; x_in <= "01100011"; z_correct<="1101101001111101";
        when 8164 => y_in <= "10011111"; x_in <= "01100100"; z_correct<="1101101000011100";
        when 8165 => y_in <= "10011111"; x_in <= "01100101"; z_correct<="1101100110111011";
        when 8166 => y_in <= "10011111"; x_in <= "01100110"; z_correct<="1101100101011010";
        when 8167 => y_in <= "10011111"; x_in <= "01100111"; z_correct<="1101100011111001";
        when 8168 => y_in <= "10011111"; x_in <= "01101000"; z_correct<="1101100010011000";
        when 8169 => y_in <= "10011111"; x_in <= "01101001"; z_correct<="1101100000110111";
        when 8170 => y_in <= "10011111"; x_in <= "01101010"; z_correct<="1101011111010110";
        when 8171 => y_in <= "10011111"; x_in <= "01101011"; z_correct<="1101011101110101";
        when 8172 => y_in <= "10011111"; x_in <= "01101100"; z_correct<="1101011100010100";
        when 8173 => y_in <= "10011111"; x_in <= "01101101"; z_correct<="1101011010110011";
        when 8174 => y_in <= "10011111"; x_in <= "01101110"; z_correct<="1101011001010010";
        when 8175 => y_in <= "10011111"; x_in <= "01101111"; z_correct<="1101010111110001";
        when 8176 => y_in <= "10011111"; x_in <= "01110000"; z_correct<="1101010110010000";
        when 8177 => y_in <= "10011111"; x_in <= "01110001"; z_correct<="1101010100101111";
        when 8178 => y_in <= "10011111"; x_in <= "01110010"; z_correct<="1101010011001110";
        when 8179 => y_in <= "10011111"; x_in <= "01110011"; z_correct<="1101010001101101";
        when 8180 => y_in <= "10011111"; x_in <= "01110100"; z_correct<="1101010000001100";
        when 8181 => y_in <= "10011111"; x_in <= "01110101"; z_correct<="1101001110101011";
        when 8182 => y_in <= "10011111"; x_in <= "01110110"; z_correct<="1101001101001010";
        when 8183 => y_in <= "10011111"; x_in <= "01110111"; z_correct<="1101001011101001";
        when 8184 => y_in <= "10011111"; x_in <= "01111000"; z_correct<="1101001010001000";
        when 8185 => y_in <= "10011111"; x_in <= "01111001"; z_correct<="1101001000100111";
        when 8186 => y_in <= "10011111"; x_in <= "01111010"; z_correct<="1101000111000110";
        when 8187 => y_in <= "10011111"; x_in <= "01111011"; z_correct<="1101000101100101";
        when 8188 => y_in <= "10011111"; x_in <= "01111100"; z_correct<="1101000100000100";
        when 8189 => y_in <= "10011111"; x_in <= "01111101"; z_correct<="1101000010100011";
        when 8190 => y_in <= "10011111"; x_in <= "01111110"; z_correct<="1101000001000010";
        when 8191 => y_in <= "10011111"; x_in <= "01111111"; z_correct<="1100111111100001";
        when 8192 => y_in <= "10100000"; x_in <= "10000000"; z_correct<="0011000000000000";
        when 8193 => y_in <= "10100000"; x_in <= "10000001"; z_correct<="0010111110100000";
        when 8194 => y_in <= "10100000"; x_in <= "10000010"; z_correct<="0010111101000000";
        when 8195 => y_in <= "10100000"; x_in <= "10000011"; z_correct<="0010111011100000";
        when 8196 => y_in <= "10100000"; x_in <= "10000100"; z_correct<="0010111010000000";
        when 8197 => y_in <= "10100000"; x_in <= "10000101"; z_correct<="0010111000100000";
        when 8198 => y_in <= "10100000"; x_in <= "10000110"; z_correct<="0010110111000000";
        when 8199 => y_in <= "10100000"; x_in <= "10000111"; z_correct<="0010110101100000";
        when 8200 => y_in <= "10100000"; x_in <= "10001000"; z_correct<="0010110100000000";
        when 8201 => y_in <= "10100000"; x_in <= "10001001"; z_correct<="0010110010100000";
        when 8202 => y_in <= "10100000"; x_in <= "10001010"; z_correct<="0010110001000000";
        when 8203 => y_in <= "10100000"; x_in <= "10001011"; z_correct<="0010101111100000";
        when 8204 => y_in <= "10100000"; x_in <= "10001100"; z_correct<="0010101110000000";
        when 8205 => y_in <= "10100000"; x_in <= "10001101"; z_correct<="0010101100100000";
        when 8206 => y_in <= "10100000"; x_in <= "10001110"; z_correct<="0010101011000000";
        when 8207 => y_in <= "10100000"; x_in <= "10001111"; z_correct<="0010101001100000";
        when 8208 => y_in <= "10100000"; x_in <= "10010000"; z_correct<="0010101000000000";
        when 8209 => y_in <= "10100000"; x_in <= "10010001"; z_correct<="0010100110100000";
        when 8210 => y_in <= "10100000"; x_in <= "10010010"; z_correct<="0010100101000000";
        when 8211 => y_in <= "10100000"; x_in <= "10010011"; z_correct<="0010100011100000";
        when 8212 => y_in <= "10100000"; x_in <= "10010100"; z_correct<="0010100010000000";
        when 8213 => y_in <= "10100000"; x_in <= "10010101"; z_correct<="0010100000100000";
        when 8214 => y_in <= "10100000"; x_in <= "10010110"; z_correct<="0010011111000000";
        when 8215 => y_in <= "10100000"; x_in <= "10010111"; z_correct<="0010011101100000";
        when 8216 => y_in <= "10100000"; x_in <= "10011000"; z_correct<="0010011100000000";
        when 8217 => y_in <= "10100000"; x_in <= "10011001"; z_correct<="0010011010100000";
        when 8218 => y_in <= "10100000"; x_in <= "10011010"; z_correct<="0010011001000000";
        when 8219 => y_in <= "10100000"; x_in <= "10011011"; z_correct<="0010010111100000";
        when 8220 => y_in <= "10100000"; x_in <= "10011100"; z_correct<="0010010110000000";
        when 8221 => y_in <= "10100000"; x_in <= "10011101"; z_correct<="0010010100100000";
        when 8222 => y_in <= "10100000"; x_in <= "10011110"; z_correct<="0010010011000000";
        when 8223 => y_in <= "10100000"; x_in <= "10011111"; z_correct<="0010010001100000";
        when 8224 => y_in <= "10100000"; x_in <= "10100000"; z_correct<="0010010000000000";
        when 8225 => y_in <= "10100000"; x_in <= "10100001"; z_correct<="0010001110100000";
        when 8226 => y_in <= "10100000"; x_in <= "10100010"; z_correct<="0010001101000000";
        when 8227 => y_in <= "10100000"; x_in <= "10100011"; z_correct<="0010001011100000";
        when 8228 => y_in <= "10100000"; x_in <= "10100100"; z_correct<="0010001010000000";
        when 8229 => y_in <= "10100000"; x_in <= "10100101"; z_correct<="0010001000100000";
        when 8230 => y_in <= "10100000"; x_in <= "10100110"; z_correct<="0010000111000000";
        when 8231 => y_in <= "10100000"; x_in <= "10100111"; z_correct<="0010000101100000";
        when 8232 => y_in <= "10100000"; x_in <= "10101000"; z_correct<="0010000100000000";
        when 8233 => y_in <= "10100000"; x_in <= "10101001"; z_correct<="0010000010100000";
        when 8234 => y_in <= "10100000"; x_in <= "10101010"; z_correct<="0010000001000000";
        when 8235 => y_in <= "10100000"; x_in <= "10101011"; z_correct<="0001111111100000";
        when 8236 => y_in <= "10100000"; x_in <= "10101100"; z_correct<="0001111110000000";
        when 8237 => y_in <= "10100000"; x_in <= "10101101"; z_correct<="0001111100100000";
        when 8238 => y_in <= "10100000"; x_in <= "10101110"; z_correct<="0001111011000000";
        when 8239 => y_in <= "10100000"; x_in <= "10101111"; z_correct<="0001111001100000";
        when 8240 => y_in <= "10100000"; x_in <= "10110000"; z_correct<="0001111000000000";
        when 8241 => y_in <= "10100000"; x_in <= "10110001"; z_correct<="0001110110100000";
        when 8242 => y_in <= "10100000"; x_in <= "10110010"; z_correct<="0001110101000000";
        when 8243 => y_in <= "10100000"; x_in <= "10110011"; z_correct<="0001110011100000";
        when 8244 => y_in <= "10100000"; x_in <= "10110100"; z_correct<="0001110010000000";
        when 8245 => y_in <= "10100000"; x_in <= "10110101"; z_correct<="0001110000100000";
        when 8246 => y_in <= "10100000"; x_in <= "10110110"; z_correct<="0001101111000000";
        when 8247 => y_in <= "10100000"; x_in <= "10110111"; z_correct<="0001101101100000";
        when 8248 => y_in <= "10100000"; x_in <= "10111000"; z_correct<="0001101100000000";
        when 8249 => y_in <= "10100000"; x_in <= "10111001"; z_correct<="0001101010100000";
        when 8250 => y_in <= "10100000"; x_in <= "10111010"; z_correct<="0001101001000000";
        when 8251 => y_in <= "10100000"; x_in <= "10111011"; z_correct<="0001100111100000";
        when 8252 => y_in <= "10100000"; x_in <= "10111100"; z_correct<="0001100110000000";
        when 8253 => y_in <= "10100000"; x_in <= "10111101"; z_correct<="0001100100100000";
        when 8254 => y_in <= "10100000"; x_in <= "10111110"; z_correct<="0001100011000000";
        when 8255 => y_in <= "10100000"; x_in <= "10111111"; z_correct<="0001100001100000";
        when 8256 => y_in <= "10100000"; x_in <= "11000000"; z_correct<="0001100000000000";
        when 8257 => y_in <= "10100000"; x_in <= "11000001"; z_correct<="0001011110100000";
        when 8258 => y_in <= "10100000"; x_in <= "11000010"; z_correct<="0001011101000000";
        when 8259 => y_in <= "10100000"; x_in <= "11000011"; z_correct<="0001011011100000";
        when 8260 => y_in <= "10100000"; x_in <= "11000100"; z_correct<="0001011010000000";
        when 8261 => y_in <= "10100000"; x_in <= "11000101"; z_correct<="0001011000100000";
        when 8262 => y_in <= "10100000"; x_in <= "11000110"; z_correct<="0001010111000000";
        when 8263 => y_in <= "10100000"; x_in <= "11000111"; z_correct<="0001010101100000";
        when 8264 => y_in <= "10100000"; x_in <= "11001000"; z_correct<="0001010100000000";
        when 8265 => y_in <= "10100000"; x_in <= "11001001"; z_correct<="0001010010100000";
        when 8266 => y_in <= "10100000"; x_in <= "11001010"; z_correct<="0001010001000000";
        when 8267 => y_in <= "10100000"; x_in <= "11001011"; z_correct<="0001001111100000";
        when 8268 => y_in <= "10100000"; x_in <= "11001100"; z_correct<="0001001110000000";
        when 8269 => y_in <= "10100000"; x_in <= "11001101"; z_correct<="0001001100100000";
        when 8270 => y_in <= "10100000"; x_in <= "11001110"; z_correct<="0001001011000000";
        when 8271 => y_in <= "10100000"; x_in <= "11001111"; z_correct<="0001001001100000";
        when 8272 => y_in <= "10100000"; x_in <= "11010000"; z_correct<="0001001000000000";
        when 8273 => y_in <= "10100000"; x_in <= "11010001"; z_correct<="0001000110100000";
        when 8274 => y_in <= "10100000"; x_in <= "11010010"; z_correct<="0001000101000000";
        when 8275 => y_in <= "10100000"; x_in <= "11010011"; z_correct<="0001000011100000";
        when 8276 => y_in <= "10100000"; x_in <= "11010100"; z_correct<="0001000010000000";
        when 8277 => y_in <= "10100000"; x_in <= "11010101"; z_correct<="0001000000100000";
        when 8278 => y_in <= "10100000"; x_in <= "11010110"; z_correct<="0000111111000000";
        when 8279 => y_in <= "10100000"; x_in <= "11010111"; z_correct<="0000111101100000";
        when 8280 => y_in <= "10100000"; x_in <= "11011000"; z_correct<="0000111100000000";
        when 8281 => y_in <= "10100000"; x_in <= "11011001"; z_correct<="0000111010100000";
        when 8282 => y_in <= "10100000"; x_in <= "11011010"; z_correct<="0000111001000000";
        when 8283 => y_in <= "10100000"; x_in <= "11011011"; z_correct<="0000110111100000";
        when 8284 => y_in <= "10100000"; x_in <= "11011100"; z_correct<="0000110110000000";
        when 8285 => y_in <= "10100000"; x_in <= "11011101"; z_correct<="0000110100100000";
        when 8286 => y_in <= "10100000"; x_in <= "11011110"; z_correct<="0000110011000000";
        when 8287 => y_in <= "10100000"; x_in <= "11011111"; z_correct<="0000110001100000";
        when 8288 => y_in <= "10100000"; x_in <= "11100000"; z_correct<="0000110000000000";
        when 8289 => y_in <= "10100000"; x_in <= "11100001"; z_correct<="0000101110100000";
        when 8290 => y_in <= "10100000"; x_in <= "11100010"; z_correct<="0000101101000000";
        when 8291 => y_in <= "10100000"; x_in <= "11100011"; z_correct<="0000101011100000";
        when 8292 => y_in <= "10100000"; x_in <= "11100100"; z_correct<="0000101010000000";
        when 8293 => y_in <= "10100000"; x_in <= "11100101"; z_correct<="0000101000100000";
        when 8294 => y_in <= "10100000"; x_in <= "11100110"; z_correct<="0000100111000000";
        when 8295 => y_in <= "10100000"; x_in <= "11100111"; z_correct<="0000100101100000";
        when 8296 => y_in <= "10100000"; x_in <= "11101000"; z_correct<="0000100100000000";
        when 8297 => y_in <= "10100000"; x_in <= "11101001"; z_correct<="0000100010100000";
        when 8298 => y_in <= "10100000"; x_in <= "11101010"; z_correct<="0000100001000000";
        when 8299 => y_in <= "10100000"; x_in <= "11101011"; z_correct<="0000011111100000";
        when 8300 => y_in <= "10100000"; x_in <= "11101100"; z_correct<="0000011110000000";
        when 8301 => y_in <= "10100000"; x_in <= "11101101"; z_correct<="0000011100100000";
        when 8302 => y_in <= "10100000"; x_in <= "11101110"; z_correct<="0000011011000000";
        when 8303 => y_in <= "10100000"; x_in <= "11101111"; z_correct<="0000011001100000";
        when 8304 => y_in <= "10100000"; x_in <= "11110000"; z_correct<="0000011000000000";
        when 8305 => y_in <= "10100000"; x_in <= "11110001"; z_correct<="0000010110100000";
        when 8306 => y_in <= "10100000"; x_in <= "11110010"; z_correct<="0000010101000000";
        when 8307 => y_in <= "10100000"; x_in <= "11110011"; z_correct<="0000010011100000";
        when 8308 => y_in <= "10100000"; x_in <= "11110100"; z_correct<="0000010010000000";
        when 8309 => y_in <= "10100000"; x_in <= "11110101"; z_correct<="0000010000100000";
        when 8310 => y_in <= "10100000"; x_in <= "11110110"; z_correct<="0000001111000000";
        when 8311 => y_in <= "10100000"; x_in <= "11110111"; z_correct<="0000001101100000";
        when 8312 => y_in <= "10100000"; x_in <= "11111000"; z_correct<="0000001100000000";
        when 8313 => y_in <= "10100000"; x_in <= "11111001"; z_correct<="0000001010100000";
        when 8314 => y_in <= "10100000"; x_in <= "11111010"; z_correct<="0000001001000000";
        when 8315 => y_in <= "10100000"; x_in <= "11111011"; z_correct<="0000000111100000";
        when 8316 => y_in <= "10100000"; x_in <= "11111100"; z_correct<="0000000110000000";
        when 8317 => y_in <= "10100000"; x_in <= "11111101"; z_correct<="0000000100100000";
        when 8318 => y_in <= "10100000"; x_in <= "11111110"; z_correct<="0000000011000000";
        when 8319 => y_in <= "10100000"; x_in <= "11111111"; z_correct<="0000000001100000";
        when 8320 => y_in <= "10100000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 8321 => y_in <= "10100000"; x_in <= "00000001"; z_correct<="1111111110100000";
        when 8322 => y_in <= "10100000"; x_in <= "00000010"; z_correct<="1111111101000000";
        when 8323 => y_in <= "10100000"; x_in <= "00000011"; z_correct<="1111111011100000";
        when 8324 => y_in <= "10100000"; x_in <= "00000100"; z_correct<="1111111010000000";
        when 8325 => y_in <= "10100000"; x_in <= "00000101"; z_correct<="1111111000100000";
        when 8326 => y_in <= "10100000"; x_in <= "00000110"; z_correct<="1111110111000000";
        when 8327 => y_in <= "10100000"; x_in <= "00000111"; z_correct<="1111110101100000";
        when 8328 => y_in <= "10100000"; x_in <= "00001000"; z_correct<="1111110100000000";
        when 8329 => y_in <= "10100000"; x_in <= "00001001"; z_correct<="1111110010100000";
        when 8330 => y_in <= "10100000"; x_in <= "00001010"; z_correct<="1111110001000000";
        when 8331 => y_in <= "10100000"; x_in <= "00001011"; z_correct<="1111101111100000";
        when 8332 => y_in <= "10100000"; x_in <= "00001100"; z_correct<="1111101110000000";
        when 8333 => y_in <= "10100000"; x_in <= "00001101"; z_correct<="1111101100100000";
        when 8334 => y_in <= "10100000"; x_in <= "00001110"; z_correct<="1111101011000000";
        when 8335 => y_in <= "10100000"; x_in <= "00001111"; z_correct<="1111101001100000";
        when 8336 => y_in <= "10100000"; x_in <= "00010000"; z_correct<="1111101000000000";
        when 8337 => y_in <= "10100000"; x_in <= "00010001"; z_correct<="1111100110100000";
        when 8338 => y_in <= "10100000"; x_in <= "00010010"; z_correct<="1111100101000000";
        when 8339 => y_in <= "10100000"; x_in <= "00010011"; z_correct<="1111100011100000";
        when 8340 => y_in <= "10100000"; x_in <= "00010100"; z_correct<="1111100010000000";
        when 8341 => y_in <= "10100000"; x_in <= "00010101"; z_correct<="1111100000100000";
        when 8342 => y_in <= "10100000"; x_in <= "00010110"; z_correct<="1111011111000000";
        when 8343 => y_in <= "10100000"; x_in <= "00010111"; z_correct<="1111011101100000";
        when 8344 => y_in <= "10100000"; x_in <= "00011000"; z_correct<="1111011100000000";
        when 8345 => y_in <= "10100000"; x_in <= "00011001"; z_correct<="1111011010100000";
        when 8346 => y_in <= "10100000"; x_in <= "00011010"; z_correct<="1111011001000000";
        when 8347 => y_in <= "10100000"; x_in <= "00011011"; z_correct<="1111010111100000";
        when 8348 => y_in <= "10100000"; x_in <= "00011100"; z_correct<="1111010110000000";
        when 8349 => y_in <= "10100000"; x_in <= "00011101"; z_correct<="1111010100100000";
        when 8350 => y_in <= "10100000"; x_in <= "00011110"; z_correct<="1111010011000000";
        when 8351 => y_in <= "10100000"; x_in <= "00011111"; z_correct<="1111010001100000";
        when 8352 => y_in <= "10100000"; x_in <= "00100000"; z_correct<="1111010000000000";
        when 8353 => y_in <= "10100000"; x_in <= "00100001"; z_correct<="1111001110100000";
        when 8354 => y_in <= "10100000"; x_in <= "00100010"; z_correct<="1111001101000000";
        when 8355 => y_in <= "10100000"; x_in <= "00100011"; z_correct<="1111001011100000";
        when 8356 => y_in <= "10100000"; x_in <= "00100100"; z_correct<="1111001010000000";
        when 8357 => y_in <= "10100000"; x_in <= "00100101"; z_correct<="1111001000100000";
        when 8358 => y_in <= "10100000"; x_in <= "00100110"; z_correct<="1111000111000000";
        when 8359 => y_in <= "10100000"; x_in <= "00100111"; z_correct<="1111000101100000";
        when 8360 => y_in <= "10100000"; x_in <= "00101000"; z_correct<="1111000100000000";
        when 8361 => y_in <= "10100000"; x_in <= "00101001"; z_correct<="1111000010100000";
        when 8362 => y_in <= "10100000"; x_in <= "00101010"; z_correct<="1111000001000000";
        when 8363 => y_in <= "10100000"; x_in <= "00101011"; z_correct<="1110111111100000";
        when 8364 => y_in <= "10100000"; x_in <= "00101100"; z_correct<="1110111110000000";
        when 8365 => y_in <= "10100000"; x_in <= "00101101"; z_correct<="1110111100100000";
        when 8366 => y_in <= "10100000"; x_in <= "00101110"; z_correct<="1110111011000000";
        when 8367 => y_in <= "10100000"; x_in <= "00101111"; z_correct<="1110111001100000";
        when 8368 => y_in <= "10100000"; x_in <= "00110000"; z_correct<="1110111000000000";
        when 8369 => y_in <= "10100000"; x_in <= "00110001"; z_correct<="1110110110100000";
        when 8370 => y_in <= "10100000"; x_in <= "00110010"; z_correct<="1110110101000000";
        when 8371 => y_in <= "10100000"; x_in <= "00110011"; z_correct<="1110110011100000";
        when 8372 => y_in <= "10100000"; x_in <= "00110100"; z_correct<="1110110010000000";
        when 8373 => y_in <= "10100000"; x_in <= "00110101"; z_correct<="1110110000100000";
        when 8374 => y_in <= "10100000"; x_in <= "00110110"; z_correct<="1110101111000000";
        when 8375 => y_in <= "10100000"; x_in <= "00110111"; z_correct<="1110101101100000";
        when 8376 => y_in <= "10100000"; x_in <= "00111000"; z_correct<="1110101100000000";
        when 8377 => y_in <= "10100000"; x_in <= "00111001"; z_correct<="1110101010100000";
        when 8378 => y_in <= "10100000"; x_in <= "00111010"; z_correct<="1110101001000000";
        when 8379 => y_in <= "10100000"; x_in <= "00111011"; z_correct<="1110100111100000";
        when 8380 => y_in <= "10100000"; x_in <= "00111100"; z_correct<="1110100110000000";
        when 8381 => y_in <= "10100000"; x_in <= "00111101"; z_correct<="1110100100100000";
        when 8382 => y_in <= "10100000"; x_in <= "00111110"; z_correct<="1110100011000000";
        when 8383 => y_in <= "10100000"; x_in <= "00111111"; z_correct<="1110100001100000";
        when 8384 => y_in <= "10100000"; x_in <= "01000000"; z_correct<="1110100000000000";
        when 8385 => y_in <= "10100000"; x_in <= "01000001"; z_correct<="1110011110100000";
        when 8386 => y_in <= "10100000"; x_in <= "01000010"; z_correct<="1110011101000000";
        when 8387 => y_in <= "10100000"; x_in <= "01000011"; z_correct<="1110011011100000";
        when 8388 => y_in <= "10100000"; x_in <= "01000100"; z_correct<="1110011010000000";
        when 8389 => y_in <= "10100000"; x_in <= "01000101"; z_correct<="1110011000100000";
        when 8390 => y_in <= "10100000"; x_in <= "01000110"; z_correct<="1110010111000000";
        when 8391 => y_in <= "10100000"; x_in <= "01000111"; z_correct<="1110010101100000";
        when 8392 => y_in <= "10100000"; x_in <= "01001000"; z_correct<="1110010100000000";
        when 8393 => y_in <= "10100000"; x_in <= "01001001"; z_correct<="1110010010100000";
        when 8394 => y_in <= "10100000"; x_in <= "01001010"; z_correct<="1110010001000000";
        when 8395 => y_in <= "10100000"; x_in <= "01001011"; z_correct<="1110001111100000";
        when 8396 => y_in <= "10100000"; x_in <= "01001100"; z_correct<="1110001110000000";
        when 8397 => y_in <= "10100000"; x_in <= "01001101"; z_correct<="1110001100100000";
        when 8398 => y_in <= "10100000"; x_in <= "01001110"; z_correct<="1110001011000000";
        when 8399 => y_in <= "10100000"; x_in <= "01001111"; z_correct<="1110001001100000";
        when 8400 => y_in <= "10100000"; x_in <= "01010000"; z_correct<="1110001000000000";
        when 8401 => y_in <= "10100000"; x_in <= "01010001"; z_correct<="1110000110100000";
        when 8402 => y_in <= "10100000"; x_in <= "01010010"; z_correct<="1110000101000000";
        when 8403 => y_in <= "10100000"; x_in <= "01010011"; z_correct<="1110000011100000";
        when 8404 => y_in <= "10100000"; x_in <= "01010100"; z_correct<="1110000010000000";
        when 8405 => y_in <= "10100000"; x_in <= "01010101"; z_correct<="1110000000100000";
        when 8406 => y_in <= "10100000"; x_in <= "01010110"; z_correct<="1101111111000000";
        when 8407 => y_in <= "10100000"; x_in <= "01010111"; z_correct<="1101111101100000";
        when 8408 => y_in <= "10100000"; x_in <= "01011000"; z_correct<="1101111100000000";
        when 8409 => y_in <= "10100000"; x_in <= "01011001"; z_correct<="1101111010100000";
        when 8410 => y_in <= "10100000"; x_in <= "01011010"; z_correct<="1101111001000000";
        when 8411 => y_in <= "10100000"; x_in <= "01011011"; z_correct<="1101110111100000";
        when 8412 => y_in <= "10100000"; x_in <= "01011100"; z_correct<="1101110110000000";
        when 8413 => y_in <= "10100000"; x_in <= "01011101"; z_correct<="1101110100100000";
        when 8414 => y_in <= "10100000"; x_in <= "01011110"; z_correct<="1101110011000000";
        when 8415 => y_in <= "10100000"; x_in <= "01011111"; z_correct<="1101110001100000";
        when 8416 => y_in <= "10100000"; x_in <= "01100000"; z_correct<="1101110000000000";
        when 8417 => y_in <= "10100000"; x_in <= "01100001"; z_correct<="1101101110100000";
        when 8418 => y_in <= "10100000"; x_in <= "01100010"; z_correct<="1101101101000000";
        when 8419 => y_in <= "10100000"; x_in <= "01100011"; z_correct<="1101101011100000";
        when 8420 => y_in <= "10100000"; x_in <= "01100100"; z_correct<="1101101010000000";
        when 8421 => y_in <= "10100000"; x_in <= "01100101"; z_correct<="1101101000100000";
        when 8422 => y_in <= "10100000"; x_in <= "01100110"; z_correct<="1101100111000000";
        when 8423 => y_in <= "10100000"; x_in <= "01100111"; z_correct<="1101100101100000";
        when 8424 => y_in <= "10100000"; x_in <= "01101000"; z_correct<="1101100100000000";
        when 8425 => y_in <= "10100000"; x_in <= "01101001"; z_correct<="1101100010100000";
        when 8426 => y_in <= "10100000"; x_in <= "01101010"; z_correct<="1101100001000000";
        when 8427 => y_in <= "10100000"; x_in <= "01101011"; z_correct<="1101011111100000";
        when 8428 => y_in <= "10100000"; x_in <= "01101100"; z_correct<="1101011110000000";
        when 8429 => y_in <= "10100000"; x_in <= "01101101"; z_correct<="1101011100100000";
        when 8430 => y_in <= "10100000"; x_in <= "01101110"; z_correct<="1101011011000000";
        when 8431 => y_in <= "10100000"; x_in <= "01101111"; z_correct<="1101011001100000";
        when 8432 => y_in <= "10100000"; x_in <= "01110000"; z_correct<="1101011000000000";
        when 8433 => y_in <= "10100000"; x_in <= "01110001"; z_correct<="1101010110100000";
        when 8434 => y_in <= "10100000"; x_in <= "01110010"; z_correct<="1101010101000000";
        when 8435 => y_in <= "10100000"; x_in <= "01110011"; z_correct<="1101010011100000";
        when 8436 => y_in <= "10100000"; x_in <= "01110100"; z_correct<="1101010010000000";
        when 8437 => y_in <= "10100000"; x_in <= "01110101"; z_correct<="1101010000100000";
        when 8438 => y_in <= "10100000"; x_in <= "01110110"; z_correct<="1101001111000000";
        when 8439 => y_in <= "10100000"; x_in <= "01110111"; z_correct<="1101001101100000";
        when 8440 => y_in <= "10100000"; x_in <= "01111000"; z_correct<="1101001100000000";
        when 8441 => y_in <= "10100000"; x_in <= "01111001"; z_correct<="1101001010100000";
        when 8442 => y_in <= "10100000"; x_in <= "01111010"; z_correct<="1101001001000000";
        when 8443 => y_in <= "10100000"; x_in <= "01111011"; z_correct<="1101000111100000";
        when 8444 => y_in <= "10100000"; x_in <= "01111100"; z_correct<="1101000110000000";
        when 8445 => y_in <= "10100000"; x_in <= "01111101"; z_correct<="1101000100100000";
        when 8446 => y_in <= "10100000"; x_in <= "01111110"; z_correct<="1101000011000000";
        when 8447 => y_in <= "10100000"; x_in <= "01111111"; z_correct<="1101000001100000";
        when 8448 => y_in <= "10100001"; x_in <= "10000000"; z_correct<="0010111110000000";
        when 8449 => y_in <= "10100001"; x_in <= "10000001"; z_correct<="0010111100100001";
        when 8450 => y_in <= "10100001"; x_in <= "10000010"; z_correct<="0010111011000010";
        when 8451 => y_in <= "10100001"; x_in <= "10000011"; z_correct<="0010111001100011";
        when 8452 => y_in <= "10100001"; x_in <= "10000100"; z_correct<="0010111000000100";
        when 8453 => y_in <= "10100001"; x_in <= "10000101"; z_correct<="0010110110100101";
        when 8454 => y_in <= "10100001"; x_in <= "10000110"; z_correct<="0010110101000110";
        when 8455 => y_in <= "10100001"; x_in <= "10000111"; z_correct<="0010110011100111";
        when 8456 => y_in <= "10100001"; x_in <= "10001000"; z_correct<="0010110010001000";
        when 8457 => y_in <= "10100001"; x_in <= "10001001"; z_correct<="0010110000101001";
        when 8458 => y_in <= "10100001"; x_in <= "10001010"; z_correct<="0010101111001010";
        when 8459 => y_in <= "10100001"; x_in <= "10001011"; z_correct<="0010101101101011";
        when 8460 => y_in <= "10100001"; x_in <= "10001100"; z_correct<="0010101100001100";
        when 8461 => y_in <= "10100001"; x_in <= "10001101"; z_correct<="0010101010101101";
        when 8462 => y_in <= "10100001"; x_in <= "10001110"; z_correct<="0010101001001110";
        when 8463 => y_in <= "10100001"; x_in <= "10001111"; z_correct<="0010100111101111";
        when 8464 => y_in <= "10100001"; x_in <= "10010000"; z_correct<="0010100110010000";
        when 8465 => y_in <= "10100001"; x_in <= "10010001"; z_correct<="0010100100110001";
        when 8466 => y_in <= "10100001"; x_in <= "10010010"; z_correct<="0010100011010010";
        when 8467 => y_in <= "10100001"; x_in <= "10010011"; z_correct<="0010100001110011";
        when 8468 => y_in <= "10100001"; x_in <= "10010100"; z_correct<="0010100000010100";
        when 8469 => y_in <= "10100001"; x_in <= "10010101"; z_correct<="0010011110110101";
        when 8470 => y_in <= "10100001"; x_in <= "10010110"; z_correct<="0010011101010110";
        when 8471 => y_in <= "10100001"; x_in <= "10010111"; z_correct<="0010011011110111";
        when 8472 => y_in <= "10100001"; x_in <= "10011000"; z_correct<="0010011010011000";
        when 8473 => y_in <= "10100001"; x_in <= "10011001"; z_correct<="0010011000111001";
        when 8474 => y_in <= "10100001"; x_in <= "10011010"; z_correct<="0010010111011010";
        when 8475 => y_in <= "10100001"; x_in <= "10011011"; z_correct<="0010010101111011";
        when 8476 => y_in <= "10100001"; x_in <= "10011100"; z_correct<="0010010100011100";
        when 8477 => y_in <= "10100001"; x_in <= "10011101"; z_correct<="0010010010111101";
        when 8478 => y_in <= "10100001"; x_in <= "10011110"; z_correct<="0010010001011110";
        when 8479 => y_in <= "10100001"; x_in <= "10011111"; z_correct<="0010001111111111";
        when 8480 => y_in <= "10100001"; x_in <= "10100000"; z_correct<="0010001110100000";
        when 8481 => y_in <= "10100001"; x_in <= "10100001"; z_correct<="0010001101000001";
        when 8482 => y_in <= "10100001"; x_in <= "10100010"; z_correct<="0010001011100010";
        when 8483 => y_in <= "10100001"; x_in <= "10100011"; z_correct<="0010001010000011";
        when 8484 => y_in <= "10100001"; x_in <= "10100100"; z_correct<="0010001000100100";
        when 8485 => y_in <= "10100001"; x_in <= "10100101"; z_correct<="0010000111000101";
        when 8486 => y_in <= "10100001"; x_in <= "10100110"; z_correct<="0010000101100110";
        when 8487 => y_in <= "10100001"; x_in <= "10100111"; z_correct<="0010000100000111";
        when 8488 => y_in <= "10100001"; x_in <= "10101000"; z_correct<="0010000010101000";
        when 8489 => y_in <= "10100001"; x_in <= "10101001"; z_correct<="0010000001001001";
        when 8490 => y_in <= "10100001"; x_in <= "10101010"; z_correct<="0001111111101010";
        when 8491 => y_in <= "10100001"; x_in <= "10101011"; z_correct<="0001111110001011";
        when 8492 => y_in <= "10100001"; x_in <= "10101100"; z_correct<="0001111100101100";
        when 8493 => y_in <= "10100001"; x_in <= "10101101"; z_correct<="0001111011001101";
        when 8494 => y_in <= "10100001"; x_in <= "10101110"; z_correct<="0001111001101110";
        when 8495 => y_in <= "10100001"; x_in <= "10101111"; z_correct<="0001111000001111";
        when 8496 => y_in <= "10100001"; x_in <= "10110000"; z_correct<="0001110110110000";
        when 8497 => y_in <= "10100001"; x_in <= "10110001"; z_correct<="0001110101010001";
        when 8498 => y_in <= "10100001"; x_in <= "10110010"; z_correct<="0001110011110010";
        when 8499 => y_in <= "10100001"; x_in <= "10110011"; z_correct<="0001110010010011";
        when 8500 => y_in <= "10100001"; x_in <= "10110100"; z_correct<="0001110000110100";
        when 8501 => y_in <= "10100001"; x_in <= "10110101"; z_correct<="0001101111010101";
        when 8502 => y_in <= "10100001"; x_in <= "10110110"; z_correct<="0001101101110110";
        when 8503 => y_in <= "10100001"; x_in <= "10110111"; z_correct<="0001101100010111";
        when 8504 => y_in <= "10100001"; x_in <= "10111000"; z_correct<="0001101010111000";
        when 8505 => y_in <= "10100001"; x_in <= "10111001"; z_correct<="0001101001011001";
        when 8506 => y_in <= "10100001"; x_in <= "10111010"; z_correct<="0001100111111010";
        when 8507 => y_in <= "10100001"; x_in <= "10111011"; z_correct<="0001100110011011";
        when 8508 => y_in <= "10100001"; x_in <= "10111100"; z_correct<="0001100100111100";
        when 8509 => y_in <= "10100001"; x_in <= "10111101"; z_correct<="0001100011011101";
        when 8510 => y_in <= "10100001"; x_in <= "10111110"; z_correct<="0001100001111110";
        when 8511 => y_in <= "10100001"; x_in <= "10111111"; z_correct<="0001100000011111";
        when 8512 => y_in <= "10100001"; x_in <= "11000000"; z_correct<="0001011111000000";
        when 8513 => y_in <= "10100001"; x_in <= "11000001"; z_correct<="0001011101100001";
        when 8514 => y_in <= "10100001"; x_in <= "11000010"; z_correct<="0001011100000010";
        when 8515 => y_in <= "10100001"; x_in <= "11000011"; z_correct<="0001011010100011";
        when 8516 => y_in <= "10100001"; x_in <= "11000100"; z_correct<="0001011001000100";
        when 8517 => y_in <= "10100001"; x_in <= "11000101"; z_correct<="0001010111100101";
        when 8518 => y_in <= "10100001"; x_in <= "11000110"; z_correct<="0001010110000110";
        when 8519 => y_in <= "10100001"; x_in <= "11000111"; z_correct<="0001010100100111";
        when 8520 => y_in <= "10100001"; x_in <= "11001000"; z_correct<="0001010011001000";
        when 8521 => y_in <= "10100001"; x_in <= "11001001"; z_correct<="0001010001101001";
        when 8522 => y_in <= "10100001"; x_in <= "11001010"; z_correct<="0001010000001010";
        when 8523 => y_in <= "10100001"; x_in <= "11001011"; z_correct<="0001001110101011";
        when 8524 => y_in <= "10100001"; x_in <= "11001100"; z_correct<="0001001101001100";
        when 8525 => y_in <= "10100001"; x_in <= "11001101"; z_correct<="0001001011101101";
        when 8526 => y_in <= "10100001"; x_in <= "11001110"; z_correct<="0001001010001110";
        when 8527 => y_in <= "10100001"; x_in <= "11001111"; z_correct<="0001001000101111";
        when 8528 => y_in <= "10100001"; x_in <= "11010000"; z_correct<="0001000111010000";
        when 8529 => y_in <= "10100001"; x_in <= "11010001"; z_correct<="0001000101110001";
        when 8530 => y_in <= "10100001"; x_in <= "11010010"; z_correct<="0001000100010010";
        when 8531 => y_in <= "10100001"; x_in <= "11010011"; z_correct<="0001000010110011";
        when 8532 => y_in <= "10100001"; x_in <= "11010100"; z_correct<="0001000001010100";
        when 8533 => y_in <= "10100001"; x_in <= "11010101"; z_correct<="0000111111110101";
        when 8534 => y_in <= "10100001"; x_in <= "11010110"; z_correct<="0000111110010110";
        when 8535 => y_in <= "10100001"; x_in <= "11010111"; z_correct<="0000111100110111";
        when 8536 => y_in <= "10100001"; x_in <= "11011000"; z_correct<="0000111011011000";
        when 8537 => y_in <= "10100001"; x_in <= "11011001"; z_correct<="0000111001111001";
        when 8538 => y_in <= "10100001"; x_in <= "11011010"; z_correct<="0000111000011010";
        when 8539 => y_in <= "10100001"; x_in <= "11011011"; z_correct<="0000110110111011";
        when 8540 => y_in <= "10100001"; x_in <= "11011100"; z_correct<="0000110101011100";
        when 8541 => y_in <= "10100001"; x_in <= "11011101"; z_correct<="0000110011111101";
        when 8542 => y_in <= "10100001"; x_in <= "11011110"; z_correct<="0000110010011110";
        when 8543 => y_in <= "10100001"; x_in <= "11011111"; z_correct<="0000110000111111";
        when 8544 => y_in <= "10100001"; x_in <= "11100000"; z_correct<="0000101111100000";
        when 8545 => y_in <= "10100001"; x_in <= "11100001"; z_correct<="0000101110000001";
        when 8546 => y_in <= "10100001"; x_in <= "11100010"; z_correct<="0000101100100010";
        when 8547 => y_in <= "10100001"; x_in <= "11100011"; z_correct<="0000101011000011";
        when 8548 => y_in <= "10100001"; x_in <= "11100100"; z_correct<="0000101001100100";
        when 8549 => y_in <= "10100001"; x_in <= "11100101"; z_correct<="0000101000000101";
        when 8550 => y_in <= "10100001"; x_in <= "11100110"; z_correct<="0000100110100110";
        when 8551 => y_in <= "10100001"; x_in <= "11100111"; z_correct<="0000100101000111";
        when 8552 => y_in <= "10100001"; x_in <= "11101000"; z_correct<="0000100011101000";
        when 8553 => y_in <= "10100001"; x_in <= "11101001"; z_correct<="0000100010001001";
        when 8554 => y_in <= "10100001"; x_in <= "11101010"; z_correct<="0000100000101010";
        when 8555 => y_in <= "10100001"; x_in <= "11101011"; z_correct<="0000011111001011";
        when 8556 => y_in <= "10100001"; x_in <= "11101100"; z_correct<="0000011101101100";
        when 8557 => y_in <= "10100001"; x_in <= "11101101"; z_correct<="0000011100001101";
        when 8558 => y_in <= "10100001"; x_in <= "11101110"; z_correct<="0000011010101110";
        when 8559 => y_in <= "10100001"; x_in <= "11101111"; z_correct<="0000011001001111";
        when 8560 => y_in <= "10100001"; x_in <= "11110000"; z_correct<="0000010111110000";
        when 8561 => y_in <= "10100001"; x_in <= "11110001"; z_correct<="0000010110010001";
        when 8562 => y_in <= "10100001"; x_in <= "11110010"; z_correct<="0000010100110010";
        when 8563 => y_in <= "10100001"; x_in <= "11110011"; z_correct<="0000010011010011";
        when 8564 => y_in <= "10100001"; x_in <= "11110100"; z_correct<="0000010001110100";
        when 8565 => y_in <= "10100001"; x_in <= "11110101"; z_correct<="0000010000010101";
        when 8566 => y_in <= "10100001"; x_in <= "11110110"; z_correct<="0000001110110110";
        when 8567 => y_in <= "10100001"; x_in <= "11110111"; z_correct<="0000001101010111";
        when 8568 => y_in <= "10100001"; x_in <= "11111000"; z_correct<="0000001011111000";
        when 8569 => y_in <= "10100001"; x_in <= "11111001"; z_correct<="0000001010011001";
        when 8570 => y_in <= "10100001"; x_in <= "11111010"; z_correct<="0000001000111010";
        when 8571 => y_in <= "10100001"; x_in <= "11111011"; z_correct<="0000000111011011";
        when 8572 => y_in <= "10100001"; x_in <= "11111100"; z_correct<="0000000101111100";
        when 8573 => y_in <= "10100001"; x_in <= "11111101"; z_correct<="0000000100011101";
        when 8574 => y_in <= "10100001"; x_in <= "11111110"; z_correct<="0000000010111110";
        when 8575 => y_in <= "10100001"; x_in <= "11111111"; z_correct<="0000000001011111";
        when 8576 => y_in <= "10100001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 8577 => y_in <= "10100001"; x_in <= "00000001"; z_correct<="1111111110100001";
        when 8578 => y_in <= "10100001"; x_in <= "00000010"; z_correct<="1111111101000010";
        when 8579 => y_in <= "10100001"; x_in <= "00000011"; z_correct<="1111111011100011";
        when 8580 => y_in <= "10100001"; x_in <= "00000100"; z_correct<="1111111010000100";
        when 8581 => y_in <= "10100001"; x_in <= "00000101"; z_correct<="1111111000100101";
        when 8582 => y_in <= "10100001"; x_in <= "00000110"; z_correct<="1111110111000110";
        when 8583 => y_in <= "10100001"; x_in <= "00000111"; z_correct<="1111110101100111";
        when 8584 => y_in <= "10100001"; x_in <= "00001000"; z_correct<="1111110100001000";
        when 8585 => y_in <= "10100001"; x_in <= "00001001"; z_correct<="1111110010101001";
        when 8586 => y_in <= "10100001"; x_in <= "00001010"; z_correct<="1111110001001010";
        when 8587 => y_in <= "10100001"; x_in <= "00001011"; z_correct<="1111101111101011";
        when 8588 => y_in <= "10100001"; x_in <= "00001100"; z_correct<="1111101110001100";
        when 8589 => y_in <= "10100001"; x_in <= "00001101"; z_correct<="1111101100101101";
        when 8590 => y_in <= "10100001"; x_in <= "00001110"; z_correct<="1111101011001110";
        when 8591 => y_in <= "10100001"; x_in <= "00001111"; z_correct<="1111101001101111";
        when 8592 => y_in <= "10100001"; x_in <= "00010000"; z_correct<="1111101000010000";
        when 8593 => y_in <= "10100001"; x_in <= "00010001"; z_correct<="1111100110110001";
        when 8594 => y_in <= "10100001"; x_in <= "00010010"; z_correct<="1111100101010010";
        when 8595 => y_in <= "10100001"; x_in <= "00010011"; z_correct<="1111100011110011";
        when 8596 => y_in <= "10100001"; x_in <= "00010100"; z_correct<="1111100010010100";
        when 8597 => y_in <= "10100001"; x_in <= "00010101"; z_correct<="1111100000110101";
        when 8598 => y_in <= "10100001"; x_in <= "00010110"; z_correct<="1111011111010110";
        when 8599 => y_in <= "10100001"; x_in <= "00010111"; z_correct<="1111011101110111";
        when 8600 => y_in <= "10100001"; x_in <= "00011000"; z_correct<="1111011100011000";
        when 8601 => y_in <= "10100001"; x_in <= "00011001"; z_correct<="1111011010111001";
        when 8602 => y_in <= "10100001"; x_in <= "00011010"; z_correct<="1111011001011010";
        when 8603 => y_in <= "10100001"; x_in <= "00011011"; z_correct<="1111010111111011";
        when 8604 => y_in <= "10100001"; x_in <= "00011100"; z_correct<="1111010110011100";
        when 8605 => y_in <= "10100001"; x_in <= "00011101"; z_correct<="1111010100111101";
        when 8606 => y_in <= "10100001"; x_in <= "00011110"; z_correct<="1111010011011110";
        when 8607 => y_in <= "10100001"; x_in <= "00011111"; z_correct<="1111010001111111";
        when 8608 => y_in <= "10100001"; x_in <= "00100000"; z_correct<="1111010000100000";
        when 8609 => y_in <= "10100001"; x_in <= "00100001"; z_correct<="1111001111000001";
        when 8610 => y_in <= "10100001"; x_in <= "00100010"; z_correct<="1111001101100010";
        when 8611 => y_in <= "10100001"; x_in <= "00100011"; z_correct<="1111001100000011";
        when 8612 => y_in <= "10100001"; x_in <= "00100100"; z_correct<="1111001010100100";
        when 8613 => y_in <= "10100001"; x_in <= "00100101"; z_correct<="1111001001000101";
        when 8614 => y_in <= "10100001"; x_in <= "00100110"; z_correct<="1111000111100110";
        when 8615 => y_in <= "10100001"; x_in <= "00100111"; z_correct<="1111000110000111";
        when 8616 => y_in <= "10100001"; x_in <= "00101000"; z_correct<="1111000100101000";
        when 8617 => y_in <= "10100001"; x_in <= "00101001"; z_correct<="1111000011001001";
        when 8618 => y_in <= "10100001"; x_in <= "00101010"; z_correct<="1111000001101010";
        when 8619 => y_in <= "10100001"; x_in <= "00101011"; z_correct<="1111000000001011";
        when 8620 => y_in <= "10100001"; x_in <= "00101100"; z_correct<="1110111110101100";
        when 8621 => y_in <= "10100001"; x_in <= "00101101"; z_correct<="1110111101001101";
        when 8622 => y_in <= "10100001"; x_in <= "00101110"; z_correct<="1110111011101110";
        when 8623 => y_in <= "10100001"; x_in <= "00101111"; z_correct<="1110111010001111";
        when 8624 => y_in <= "10100001"; x_in <= "00110000"; z_correct<="1110111000110000";
        when 8625 => y_in <= "10100001"; x_in <= "00110001"; z_correct<="1110110111010001";
        when 8626 => y_in <= "10100001"; x_in <= "00110010"; z_correct<="1110110101110010";
        when 8627 => y_in <= "10100001"; x_in <= "00110011"; z_correct<="1110110100010011";
        when 8628 => y_in <= "10100001"; x_in <= "00110100"; z_correct<="1110110010110100";
        when 8629 => y_in <= "10100001"; x_in <= "00110101"; z_correct<="1110110001010101";
        when 8630 => y_in <= "10100001"; x_in <= "00110110"; z_correct<="1110101111110110";
        when 8631 => y_in <= "10100001"; x_in <= "00110111"; z_correct<="1110101110010111";
        when 8632 => y_in <= "10100001"; x_in <= "00111000"; z_correct<="1110101100111000";
        when 8633 => y_in <= "10100001"; x_in <= "00111001"; z_correct<="1110101011011001";
        when 8634 => y_in <= "10100001"; x_in <= "00111010"; z_correct<="1110101001111010";
        when 8635 => y_in <= "10100001"; x_in <= "00111011"; z_correct<="1110101000011011";
        when 8636 => y_in <= "10100001"; x_in <= "00111100"; z_correct<="1110100110111100";
        when 8637 => y_in <= "10100001"; x_in <= "00111101"; z_correct<="1110100101011101";
        when 8638 => y_in <= "10100001"; x_in <= "00111110"; z_correct<="1110100011111110";
        when 8639 => y_in <= "10100001"; x_in <= "00111111"; z_correct<="1110100010011111";
        when 8640 => y_in <= "10100001"; x_in <= "01000000"; z_correct<="1110100001000000";
        when 8641 => y_in <= "10100001"; x_in <= "01000001"; z_correct<="1110011111100001";
        when 8642 => y_in <= "10100001"; x_in <= "01000010"; z_correct<="1110011110000010";
        when 8643 => y_in <= "10100001"; x_in <= "01000011"; z_correct<="1110011100100011";
        when 8644 => y_in <= "10100001"; x_in <= "01000100"; z_correct<="1110011011000100";
        when 8645 => y_in <= "10100001"; x_in <= "01000101"; z_correct<="1110011001100101";
        when 8646 => y_in <= "10100001"; x_in <= "01000110"; z_correct<="1110011000000110";
        when 8647 => y_in <= "10100001"; x_in <= "01000111"; z_correct<="1110010110100111";
        when 8648 => y_in <= "10100001"; x_in <= "01001000"; z_correct<="1110010101001000";
        when 8649 => y_in <= "10100001"; x_in <= "01001001"; z_correct<="1110010011101001";
        when 8650 => y_in <= "10100001"; x_in <= "01001010"; z_correct<="1110010010001010";
        when 8651 => y_in <= "10100001"; x_in <= "01001011"; z_correct<="1110010000101011";
        when 8652 => y_in <= "10100001"; x_in <= "01001100"; z_correct<="1110001111001100";
        when 8653 => y_in <= "10100001"; x_in <= "01001101"; z_correct<="1110001101101101";
        when 8654 => y_in <= "10100001"; x_in <= "01001110"; z_correct<="1110001100001110";
        when 8655 => y_in <= "10100001"; x_in <= "01001111"; z_correct<="1110001010101111";
        when 8656 => y_in <= "10100001"; x_in <= "01010000"; z_correct<="1110001001010000";
        when 8657 => y_in <= "10100001"; x_in <= "01010001"; z_correct<="1110000111110001";
        when 8658 => y_in <= "10100001"; x_in <= "01010010"; z_correct<="1110000110010010";
        when 8659 => y_in <= "10100001"; x_in <= "01010011"; z_correct<="1110000100110011";
        when 8660 => y_in <= "10100001"; x_in <= "01010100"; z_correct<="1110000011010100";
        when 8661 => y_in <= "10100001"; x_in <= "01010101"; z_correct<="1110000001110101";
        when 8662 => y_in <= "10100001"; x_in <= "01010110"; z_correct<="1110000000010110";
        when 8663 => y_in <= "10100001"; x_in <= "01010111"; z_correct<="1101111110110111";
        when 8664 => y_in <= "10100001"; x_in <= "01011000"; z_correct<="1101111101011000";
        when 8665 => y_in <= "10100001"; x_in <= "01011001"; z_correct<="1101111011111001";
        when 8666 => y_in <= "10100001"; x_in <= "01011010"; z_correct<="1101111010011010";
        when 8667 => y_in <= "10100001"; x_in <= "01011011"; z_correct<="1101111000111011";
        when 8668 => y_in <= "10100001"; x_in <= "01011100"; z_correct<="1101110111011100";
        when 8669 => y_in <= "10100001"; x_in <= "01011101"; z_correct<="1101110101111101";
        when 8670 => y_in <= "10100001"; x_in <= "01011110"; z_correct<="1101110100011110";
        when 8671 => y_in <= "10100001"; x_in <= "01011111"; z_correct<="1101110010111111";
        when 8672 => y_in <= "10100001"; x_in <= "01100000"; z_correct<="1101110001100000";
        when 8673 => y_in <= "10100001"; x_in <= "01100001"; z_correct<="1101110000000001";
        when 8674 => y_in <= "10100001"; x_in <= "01100010"; z_correct<="1101101110100010";
        when 8675 => y_in <= "10100001"; x_in <= "01100011"; z_correct<="1101101101000011";
        when 8676 => y_in <= "10100001"; x_in <= "01100100"; z_correct<="1101101011100100";
        when 8677 => y_in <= "10100001"; x_in <= "01100101"; z_correct<="1101101010000101";
        when 8678 => y_in <= "10100001"; x_in <= "01100110"; z_correct<="1101101000100110";
        when 8679 => y_in <= "10100001"; x_in <= "01100111"; z_correct<="1101100111000111";
        when 8680 => y_in <= "10100001"; x_in <= "01101000"; z_correct<="1101100101101000";
        when 8681 => y_in <= "10100001"; x_in <= "01101001"; z_correct<="1101100100001001";
        when 8682 => y_in <= "10100001"; x_in <= "01101010"; z_correct<="1101100010101010";
        when 8683 => y_in <= "10100001"; x_in <= "01101011"; z_correct<="1101100001001011";
        when 8684 => y_in <= "10100001"; x_in <= "01101100"; z_correct<="1101011111101100";
        when 8685 => y_in <= "10100001"; x_in <= "01101101"; z_correct<="1101011110001101";
        when 8686 => y_in <= "10100001"; x_in <= "01101110"; z_correct<="1101011100101110";
        when 8687 => y_in <= "10100001"; x_in <= "01101111"; z_correct<="1101011011001111";
        when 8688 => y_in <= "10100001"; x_in <= "01110000"; z_correct<="1101011001110000";
        when 8689 => y_in <= "10100001"; x_in <= "01110001"; z_correct<="1101011000010001";
        when 8690 => y_in <= "10100001"; x_in <= "01110010"; z_correct<="1101010110110010";
        when 8691 => y_in <= "10100001"; x_in <= "01110011"; z_correct<="1101010101010011";
        when 8692 => y_in <= "10100001"; x_in <= "01110100"; z_correct<="1101010011110100";
        when 8693 => y_in <= "10100001"; x_in <= "01110101"; z_correct<="1101010010010101";
        when 8694 => y_in <= "10100001"; x_in <= "01110110"; z_correct<="1101010000110110";
        when 8695 => y_in <= "10100001"; x_in <= "01110111"; z_correct<="1101001111010111";
        when 8696 => y_in <= "10100001"; x_in <= "01111000"; z_correct<="1101001101111000";
        when 8697 => y_in <= "10100001"; x_in <= "01111001"; z_correct<="1101001100011001";
        when 8698 => y_in <= "10100001"; x_in <= "01111010"; z_correct<="1101001010111010";
        when 8699 => y_in <= "10100001"; x_in <= "01111011"; z_correct<="1101001001011011";
        when 8700 => y_in <= "10100001"; x_in <= "01111100"; z_correct<="1101000111111100";
        when 8701 => y_in <= "10100001"; x_in <= "01111101"; z_correct<="1101000110011101";
        when 8702 => y_in <= "10100001"; x_in <= "01111110"; z_correct<="1101000100111110";
        when 8703 => y_in <= "10100001"; x_in <= "01111111"; z_correct<="1101000011011111";
        when 8704 => y_in <= "10100010"; x_in <= "10000000"; z_correct<="0010111100000000";
        when 8705 => y_in <= "10100010"; x_in <= "10000001"; z_correct<="0010111010100010";
        when 8706 => y_in <= "10100010"; x_in <= "10000010"; z_correct<="0010111001000100";
        when 8707 => y_in <= "10100010"; x_in <= "10000011"; z_correct<="0010110111100110";
        when 8708 => y_in <= "10100010"; x_in <= "10000100"; z_correct<="0010110110001000";
        when 8709 => y_in <= "10100010"; x_in <= "10000101"; z_correct<="0010110100101010";
        when 8710 => y_in <= "10100010"; x_in <= "10000110"; z_correct<="0010110011001100";
        when 8711 => y_in <= "10100010"; x_in <= "10000111"; z_correct<="0010110001101110";
        when 8712 => y_in <= "10100010"; x_in <= "10001000"; z_correct<="0010110000010000";
        when 8713 => y_in <= "10100010"; x_in <= "10001001"; z_correct<="0010101110110010";
        when 8714 => y_in <= "10100010"; x_in <= "10001010"; z_correct<="0010101101010100";
        when 8715 => y_in <= "10100010"; x_in <= "10001011"; z_correct<="0010101011110110";
        when 8716 => y_in <= "10100010"; x_in <= "10001100"; z_correct<="0010101010011000";
        when 8717 => y_in <= "10100010"; x_in <= "10001101"; z_correct<="0010101000111010";
        when 8718 => y_in <= "10100010"; x_in <= "10001110"; z_correct<="0010100111011100";
        when 8719 => y_in <= "10100010"; x_in <= "10001111"; z_correct<="0010100101111110";
        when 8720 => y_in <= "10100010"; x_in <= "10010000"; z_correct<="0010100100100000";
        when 8721 => y_in <= "10100010"; x_in <= "10010001"; z_correct<="0010100011000010";
        when 8722 => y_in <= "10100010"; x_in <= "10010010"; z_correct<="0010100001100100";
        when 8723 => y_in <= "10100010"; x_in <= "10010011"; z_correct<="0010100000000110";
        when 8724 => y_in <= "10100010"; x_in <= "10010100"; z_correct<="0010011110101000";
        when 8725 => y_in <= "10100010"; x_in <= "10010101"; z_correct<="0010011101001010";
        when 8726 => y_in <= "10100010"; x_in <= "10010110"; z_correct<="0010011011101100";
        when 8727 => y_in <= "10100010"; x_in <= "10010111"; z_correct<="0010011010001110";
        when 8728 => y_in <= "10100010"; x_in <= "10011000"; z_correct<="0010011000110000";
        when 8729 => y_in <= "10100010"; x_in <= "10011001"; z_correct<="0010010111010010";
        when 8730 => y_in <= "10100010"; x_in <= "10011010"; z_correct<="0010010101110100";
        when 8731 => y_in <= "10100010"; x_in <= "10011011"; z_correct<="0010010100010110";
        when 8732 => y_in <= "10100010"; x_in <= "10011100"; z_correct<="0010010010111000";
        when 8733 => y_in <= "10100010"; x_in <= "10011101"; z_correct<="0010010001011010";
        when 8734 => y_in <= "10100010"; x_in <= "10011110"; z_correct<="0010001111111100";
        when 8735 => y_in <= "10100010"; x_in <= "10011111"; z_correct<="0010001110011110";
        when 8736 => y_in <= "10100010"; x_in <= "10100000"; z_correct<="0010001101000000";
        when 8737 => y_in <= "10100010"; x_in <= "10100001"; z_correct<="0010001011100010";
        when 8738 => y_in <= "10100010"; x_in <= "10100010"; z_correct<="0010001010000100";
        when 8739 => y_in <= "10100010"; x_in <= "10100011"; z_correct<="0010001000100110";
        when 8740 => y_in <= "10100010"; x_in <= "10100100"; z_correct<="0010000111001000";
        when 8741 => y_in <= "10100010"; x_in <= "10100101"; z_correct<="0010000101101010";
        when 8742 => y_in <= "10100010"; x_in <= "10100110"; z_correct<="0010000100001100";
        when 8743 => y_in <= "10100010"; x_in <= "10100111"; z_correct<="0010000010101110";
        when 8744 => y_in <= "10100010"; x_in <= "10101000"; z_correct<="0010000001010000";
        when 8745 => y_in <= "10100010"; x_in <= "10101001"; z_correct<="0001111111110010";
        when 8746 => y_in <= "10100010"; x_in <= "10101010"; z_correct<="0001111110010100";
        when 8747 => y_in <= "10100010"; x_in <= "10101011"; z_correct<="0001111100110110";
        when 8748 => y_in <= "10100010"; x_in <= "10101100"; z_correct<="0001111011011000";
        when 8749 => y_in <= "10100010"; x_in <= "10101101"; z_correct<="0001111001111010";
        when 8750 => y_in <= "10100010"; x_in <= "10101110"; z_correct<="0001111000011100";
        when 8751 => y_in <= "10100010"; x_in <= "10101111"; z_correct<="0001110110111110";
        when 8752 => y_in <= "10100010"; x_in <= "10110000"; z_correct<="0001110101100000";
        when 8753 => y_in <= "10100010"; x_in <= "10110001"; z_correct<="0001110100000010";
        when 8754 => y_in <= "10100010"; x_in <= "10110010"; z_correct<="0001110010100100";
        when 8755 => y_in <= "10100010"; x_in <= "10110011"; z_correct<="0001110001000110";
        when 8756 => y_in <= "10100010"; x_in <= "10110100"; z_correct<="0001101111101000";
        when 8757 => y_in <= "10100010"; x_in <= "10110101"; z_correct<="0001101110001010";
        when 8758 => y_in <= "10100010"; x_in <= "10110110"; z_correct<="0001101100101100";
        when 8759 => y_in <= "10100010"; x_in <= "10110111"; z_correct<="0001101011001110";
        when 8760 => y_in <= "10100010"; x_in <= "10111000"; z_correct<="0001101001110000";
        when 8761 => y_in <= "10100010"; x_in <= "10111001"; z_correct<="0001101000010010";
        when 8762 => y_in <= "10100010"; x_in <= "10111010"; z_correct<="0001100110110100";
        when 8763 => y_in <= "10100010"; x_in <= "10111011"; z_correct<="0001100101010110";
        when 8764 => y_in <= "10100010"; x_in <= "10111100"; z_correct<="0001100011111000";
        when 8765 => y_in <= "10100010"; x_in <= "10111101"; z_correct<="0001100010011010";
        when 8766 => y_in <= "10100010"; x_in <= "10111110"; z_correct<="0001100000111100";
        when 8767 => y_in <= "10100010"; x_in <= "10111111"; z_correct<="0001011111011110";
        when 8768 => y_in <= "10100010"; x_in <= "11000000"; z_correct<="0001011110000000";
        when 8769 => y_in <= "10100010"; x_in <= "11000001"; z_correct<="0001011100100010";
        when 8770 => y_in <= "10100010"; x_in <= "11000010"; z_correct<="0001011011000100";
        when 8771 => y_in <= "10100010"; x_in <= "11000011"; z_correct<="0001011001100110";
        when 8772 => y_in <= "10100010"; x_in <= "11000100"; z_correct<="0001011000001000";
        when 8773 => y_in <= "10100010"; x_in <= "11000101"; z_correct<="0001010110101010";
        when 8774 => y_in <= "10100010"; x_in <= "11000110"; z_correct<="0001010101001100";
        when 8775 => y_in <= "10100010"; x_in <= "11000111"; z_correct<="0001010011101110";
        when 8776 => y_in <= "10100010"; x_in <= "11001000"; z_correct<="0001010010010000";
        when 8777 => y_in <= "10100010"; x_in <= "11001001"; z_correct<="0001010000110010";
        when 8778 => y_in <= "10100010"; x_in <= "11001010"; z_correct<="0001001111010100";
        when 8779 => y_in <= "10100010"; x_in <= "11001011"; z_correct<="0001001101110110";
        when 8780 => y_in <= "10100010"; x_in <= "11001100"; z_correct<="0001001100011000";
        when 8781 => y_in <= "10100010"; x_in <= "11001101"; z_correct<="0001001010111010";
        when 8782 => y_in <= "10100010"; x_in <= "11001110"; z_correct<="0001001001011100";
        when 8783 => y_in <= "10100010"; x_in <= "11001111"; z_correct<="0001000111111110";
        when 8784 => y_in <= "10100010"; x_in <= "11010000"; z_correct<="0001000110100000";
        when 8785 => y_in <= "10100010"; x_in <= "11010001"; z_correct<="0001000101000010";
        when 8786 => y_in <= "10100010"; x_in <= "11010010"; z_correct<="0001000011100100";
        when 8787 => y_in <= "10100010"; x_in <= "11010011"; z_correct<="0001000010000110";
        when 8788 => y_in <= "10100010"; x_in <= "11010100"; z_correct<="0001000000101000";
        when 8789 => y_in <= "10100010"; x_in <= "11010101"; z_correct<="0000111111001010";
        when 8790 => y_in <= "10100010"; x_in <= "11010110"; z_correct<="0000111101101100";
        when 8791 => y_in <= "10100010"; x_in <= "11010111"; z_correct<="0000111100001110";
        when 8792 => y_in <= "10100010"; x_in <= "11011000"; z_correct<="0000111010110000";
        when 8793 => y_in <= "10100010"; x_in <= "11011001"; z_correct<="0000111001010010";
        when 8794 => y_in <= "10100010"; x_in <= "11011010"; z_correct<="0000110111110100";
        when 8795 => y_in <= "10100010"; x_in <= "11011011"; z_correct<="0000110110010110";
        when 8796 => y_in <= "10100010"; x_in <= "11011100"; z_correct<="0000110100111000";
        when 8797 => y_in <= "10100010"; x_in <= "11011101"; z_correct<="0000110011011010";
        when 8798 => y_in <= "10100010"; x_in <= "11011110"; z_correct<="0000110001111100";
        when 8799 => y_in <= "10100010"; x_in <= "11011111"; z_correct<="0000110000011110";
        when 8800 => y_in <= "10100010"; x_in <= "11100000"; z_correct<="0000101111000000";
        when 8801 => y_in <= "10100010"; x_in <= "11100001"; z_correct<="0000101101100010";
        when 8802 => y_in <= "10100010"; x_in <= "11100010"; z_correct<="0000101100000100";
        when 8803 => y_in <= "10100010"; x_in <= "11100011"; z_correct<="0000101010100110";
        when 8804 => y_in <= "10100010"; x_in <= "11100100"; z_correct<="0000101001001000";
        when 8805 => y_in <= "10100010"; x_in <= "11100101"; z_correct<="0000100111101010";
        when 8806 => y_in <= "10100010"; x_in <= "11100110"; z_correct<="0000100110001100";
        when 8807 => y_in <= "10100010"; x_in <= "11100111"; z_correct<="0000100100101110";
        when 8808 => y_in <= "10100010"; x_in <= "11101000"; z_correct<="0000100011010000";
        when 8809 => y_in <= "10100010"; x_in <= "11101001"; z_correct<="0000100001110010";
        when 8810 => y_in <= "10100010"; x_in <= "11101010"; z_correct<="0000100000010100";
        when 8811 => y_in <= "10100010"; x_in <= "11101011"; z_correct<="0000011110110110";
        when 8812 => y_in <= "10100010"; x_in <= "11101100"; z_correct<="0000011101011000";
        when 8813 => y_in <= "10100010"; x_in <= "11101101"; z_correct<="0000011011111010";
        when 8814 => y_in <= "10100010"; x_in <= "11101110"; z_correct<="0000011010011100";
        when 8815 => y_in <= "10100010"; x_in <= "11101111"; z_correct<="0000011000111110";
        when 8816 => y_in <= "10100010"; x_in <= "11110000"; z_correct<="0000010111100000";
        when 8817 => y_in <= "10100010"; x_in <= "11110001"; z_correct<="0000010110000010";
        when 8818 => y_in <= "10100010"; x_in <= "11110010"; z_correct<="0000010100100100";
        when 8819 => y_in <= "10100010"; x_in <= "11110011"; z_correct<="0000010011000110";
        when 8820 => y_in <= "10100010"; x_in <= "11110100"; z_correct<="0000010001101000";
        when 8821 => y_in <= "10100010"; x_in <= "11110101"; z_correct<="0000010000001010";
        when 8822 => y_in <= "10100010"; x_in <= "11110110"; z_correct<="0000001110101100";
        when 8823 => y_in <= "10100010"; x_in <= "11110111"; z_correct<="0000001101001110";
        when 8824 => y_in <= "10100010"; x_in <= "11111000"; z_correct<="0000001011110000";
        when 8825 => y_in <= "10100010"; x_in <= "11111001"; z_correct<="0000001010010010";
        when 8826 => y_in <= "10100010"; x_in <= "11111010"; z_correct<="0000001000110100";
        when 8827 => y_in <= "10100010"; x_in <= "11111011"; z_correct<="0000000111010110";
        when 8828 => y_in <= "10100010"; x_in <= "11111100"; z_correct<="0000000101111000";
        when 8829 => y_in <= "10100010"; x_in <= "11111101"; z_correct<="0000000100011010";
        when 8830 => y_in <= "10100010"; x_in <= "11111110"; z_correct<="0000000010111100";
        when 8831 => y_in <= "10100010"; x_in <= "11111111"; z_correct<="0000000001011110";
        when 8832 => y_in <= "10100010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 8833 => y_in <= "10100010"; x_in <= "00000001"; z_correct<="1111111110100010";
        when 8834 => y_in <= "10100010"; x_in <= "00000010"; z_correct<="1111111101000100";
        when 8835 => y_in <= "10100010"; x_in <= "00000011"; z_correct<="1111111011100110";
        when 8836 => y_in <= "10100010"; x_in <= "00000100"; z_correct<="1111111010001000";
        when 8837 => y_in <= "10100010"; x_in <= "00000101"; z_correct<="1111111000101010";
        when 8838 => y_in <= "10100010"; x_in <= "00000110"; z_correct<="1111110111001100";
        when 8839 => y_in <= "10100010"; x_in <= "00000111"; z_correct<="1111110101101110";
        when 8840 => y_in <= "10100010"; x_in <= "00001000"; z_correct<="1111110100010000";
        when 8841 => y_in <= "10100010"; x_in <= "00001001"; z_correct<="1111110010110010";
        when 8842 => y_in <= "10100010"; x_in <= "00001010"; z_correct<="1111110001010100";
        when 8843 => y_in <= "10100010"; x_in <= "00001011"; z_correct<="1111101111110110";
        when 8844 => y_in <= "10100010"; x_in <= "00001100"; z_correct<="1111101110011000";
        when 8845 => y_in <= "10100010"; x_in <= "00001101"; z_correct<="1111101100111010";
        when 8846 => y_in <= "10100010"; x_in <= "00001110"; z_correct<="1111101011011100";
        when 8847 => y_in <= "10100010"; x_in <= "00001111"; z_correct<="1111101001111110";
        when 8848 => y_in <= "10100010"; x_in <= "00010000"; z_correct<="1111101000100000";
        when 8849 => y_in <= "10100010"; x_in <= "00010001"; z_correct<="1111100111000010";
        when 8850 => y_in <= "10100010"; x_in <= "00010010"; z_correct<="1111100101100100";
        when 8851 => y_in <= "10100010"; x_in <= "00010011"; z_correct<="1111100100000110";
        when 8852 => y_in <= "10100010"; x_in <= "00010100"; z_correct<="1111100010101000";
        when 8853 => y_in <= "10100010"; x_in <= "00010101"; z_correct<="1111100001001010";
        when 8854 => y_in <= "10100010"; x_in <= "00010110"; z_correct<="1111011111101100";
        when 8855 => y_in <= "10100010"; x_in <= "00010111"; z_correct<="1111011110001110";
        when 8856 => y_in <= "10100010"; x_in <= "00011000"; z_correct<="1111011100110000";
        when 8857 => y_in <= "10100010"; x_in <= "00011001"; z_correct<="1111011011010010";
        when 8858 => y_in <= "10100010"; x_in <= "00011010"; z_correct<="1111011001110100";
        when 8859 => y_in <= "10100010"; x_in <= "00011011"; z_correct<="1111011000010110";
        when 8860 => y_in <= "10100010"; x_in <= "00011100"; z_correct<="1111010110111000";
        when 8861 => y_in <= "10100010"; x_in <= "00011101"; z_correct<="1111010101011010";
        when 8862 => y_in <= "10100010"; x_in <= "00011110"; z_correct<="1111010011111100";
        when 8863 => y_in <= "10100010"; x_in <= "00011111"; z_correct<="1111010010011110";
        when 8864 => y_in <= "10100010"; x_in <= "00100000"; z_correct<="1111010001000000";
        when 8865 => y_in <= "10100010"; x_in <= "00100001"; z_correct<="1111001111100010";
        when 8866 => y_in <= "10100010"; x_in <= "00100010"; z_correct<="1111001110000100";
        when 8867 => y_in <= "10100010"; x_in <= "00100011"; z_correct<="1111001100100110";
        when 8868 => y_in <= "10100010"; x_in <= "00100100"; z_correct<="1111001011001000";
        when 8869 => y_in <= "10100010"; x_in <= "00100101"; z_correct<="1111001001101010";
        when 8870 => y_in <= "10100010"; x_in <= "00100110"; z_correct<="1111001000001100";
        when 8871 => y_in <= "10100010"; x_in <= "00100111"; z_correct<="1111000110101110";
        when 8872 => y_in <= "10100010"; x_in <= "00101000"; z_correct<="1111000101010000";
        when 8873 => y_in <= "10100010"; x_in <= "00101001"; z_correct<="1111000011110010";
        when 8874 => y_in <= "10100010"; x_in <= "00101010"; z_correct<="1111000010010100";
        when 8875 => y_in <= "10100010"; x_in <= "00101011"; z_correct<="1111000000110110";
        when 8876 => y_in <= "10100010"; x_in <= "00101100"; z_correct<="1110111111011000";
        when 8877 => y_in <= "10100010"; x_in <= "00101101"; z_correct<="1110111101111010";
        when 8878 => y_in <= "10100010"; x_in <= "00101110"; z_correct<="1110111100011100";
        when 8879 => y_in <= "10100010"; x_in <= "00101111"; z_correct<="1110111010111110";
        when 8880 => y_in <= "10100010"; x_in <= "00110000"; z_correct<="1110111001100000";
        when 8881 => y_in <= "10100010"; x_in <= "00110001"; z_correct<="1110111000000010";
        when 8882 => y_in <= "10100010"; x_in <= "00110010"; z_correct<="1110110110100100";
        when 8883 => y_in <= "10100010"; x_in <= "00110011"; z_correct<="1110110101000110";
        when 8884 => y_in <= "10100010"; x_in <= "00110100"; z_correct<="1110110011101000";
        when 8885 => y_in <= "10100010"; x_in <= "00110101"; z_correct<="1110110010001010";
        when 8886 => y_in <= "10100010"; x_in <= "00110110"; z_correct<="1110110000101100";
        when 8887 => y_in <= "10100010"; x_in <= "00110111"; z_correct<="1110101111001110";
        when 8888 => y_in <= "10100010"; x_in <= "00111000"; z_correct<="1110101101110000";
        when 8889 => y_in <= "10100010"; x_in <= "00111001"; z_correct<="1110101100010010";
        when 8890 => y_in <= "10100010"; x_in <= "00111010"; z_correct<="1110101010110100";
        when 8891 => y_in <= "10100010"; x_in <= "00111011"; z_correct<="1110101001010110";
        when 8892 => y_in <= "10100010"; x_in <= "00111100"; z_correct<="1110100111111000";
        when 8893 => y_in <= "10100010"; x_in <= "00111101"; z_correct<="1110100110011010";
        when 8894 => y_in <= "10100010"; x_in <= "00111110"; z_correct<="1110100100111100";
        when 8895 => y_in <= "10100010"; x_in <= "00111111"; z_correct<="1110100011011110";
        when 8896 => y_in <= "10100010"; x_in <= "01000000"; z_correct<="1110100010000000";
        when 8897 => y_in <= "10100010"; x_in <= "01000001"; z_correct<="1110100000100010";
        when 8898 => y_in <= "10100010"; x_in <= "01000010"; z_correct<="1110011111000100";
        when 8899 => y_in <= "10100010"; x_in <= "01000011"; z_correct<="1110011101100110";
        when 8900 => y_in <= "10100010"; x_in <= "01000100"; z_correct<="1110011100001000";
        when 8901 => y_in <= "10100010"; x_in <= "01000101"; z_correct<="1110011010101010";
        when 8902 => y_in <= "10100010"; x_in <= "01000110"; z_correct<="1110011001001100";
        when 8903 => y_in <= "10100010"; x_in <= "01000111"; z_correct<="1110010111101110";
        when 8904 => y_in <= "10100010"; x_in <= "01001000"; z_correct<="1110010110010000";
        when 8905 => y_in <= "10100010"; x_in <= "01001001"; z_correct<="1110010100110010";
        when 8906 => y_in <= "10100010"; x_in <= "01001010"; z_correct<="1110010011010100";
        when 8907 => y_in <= "10100010"; x_in <= "01001011"; z_correct<="1110010001110110";
        when 8908 => y_in <= "10100010"; x_in <= "01001100"; z_correct<="1110010000011000";
        when 8909 => y_in <= "10100010"; x_in <= "01001101"; z_correct<="1110001110111010";
        when 8910 => y_in <= "10100010"; x_in <= "01001110"; z_correct<="1110001101011100";
        when 8911 => y_in <= "10100010"; x_in <= "01001111"; z_correct<="1110001011111110";
        when 8912 => y_in <= "10100010"; x_in <= "01010000"; z_correct<="1110001010100000";
        when 8913 => y_in <= "10100010"; x_in <= "01010001"; z_correct<="1110001001000010";
        when 8914 => y_in <= "10100010"; x_in <= "01010010"; z_correct<="1110000111100100";
        when 8915 => y_in <= "10100010"; x_in <= "01010011"; z_correct<="1110000110000110";
        when 8916 => y_in <= "10100010"; x_in <= "01010100"; z_correct<="1110000100101000";
        when 8917 => y_in <= "10100010"; x_in <= "01010101"; z_correct<="1110000011001010";
        when 8918 => y_in <= "10100010"; x_in <= "01010110"; z_correct<="1110000001101100";
        when 8919 => y_in <= "10100010"; x_in <= "01010111"; z_correct<="1110000000001110";
        when 8920 => y_in <= "10100010"; x_in <= "01011000"; z_correct<="1101111110110000";
        when 8921 => y_in <= "10100010"; x_in <= "01011001"; z_correct<="1101111101010010";
        when 8922 => y_in <= "10100010"; x_in <= "01011010"; z_correct<="1101111011110100";
        when 8923 => y_in <= "10100010"; x_in <= "01011011"; z_correct<="1101111010010110";
        when 8924 => y_in <= "10100010"; x_in <= "01011100"; z_correct<="1101111000111000";
        when 8925 => y_in <= "10100010"; x_in <= "01011101"; z_correct<="1101110111011010";
        when 8926 => y_in <= "10100010"; x_in <= "01011110"; z_correct<="1101110101111100";
        when 8927 => y_in <= "10100010"; x_in <= "01011111"; z_correct<="1101110100011110";
        when 8928 => y_in <= "10100010"; x_in <= "01100000"; z_correct<="1101110011000000";
        when 8929 => y_in <= "10100010"; x_in <= "01100001"; z_correct<="1101110001100010";
        when 8930 => y_in <= "10100010"; x_in <= "01100010"; z_correct<="1101110000000100";
        when 8931 => y_in <= "10100010"; x_in <= "01100011"; z_correct<="1101101110100110";
        when 8932 => y_in <= "10100010"; x_in <= "01100100"; z_correct<="1101101101001000";
        when 8933 => y_in <= "10100010"; x_in <= "01100101"; z_correct<="1101101011101010";
        when 8934 => y_in <= "10100010"; x_in <= "01100110"; z_correct<="1101101010001100";
        when 8935 => y_in <= "10100010"; x_in <= "01100111"; z_correct<="1101101000101110";
        when 8936 => y_in <= "10100010"; x_in <= "01101000"; z_correct<="1101100111010000";
        when 8937 => y_in <= "10100010"; x_in <= "01101001"; z_correct<="1101100101110010";
        when 8938 => y_in <= "10100010"; x_in <= "01101010"; z_correct<="1101100100010100";
        when 8939 => y_in <= "10100010"; x_in <= "01101011"; z_correct<="1101100010110110";
        when 8940 => y_in <= "10100010"; x_in <= "01101100"; z_correct<="1101100001011000";
        when 8941 => y_in <= "10100010"; x_in <= "01101101"; z_correct<="1101011111111010";
        when 8942 => y_in <= "10100010"; x_in <= "01101110"; z_correct<="1101011110011100";
        when 8943 => y_in <= "10100010"; x_in <= "01101111"; z_correct<="1101011100111110";
        when 8944 => y_in <= "10100010"; x_in <= "01110000"; z_correct<="1101011011100000";
        when 8945 => y_in <= "10100010"; x_in <= "01110001"; z_correct<="1101011010000010";
        when 8946 => y_in <= "10100010"; x_in <= "01110010"; z_correct<="1101011000100100";
        when 8947 => y_in <= "10100010"; x_in <= "01110011"; z_correct<="1101010111000110";
        when 8948 => y_in <= "10100010"; x_in <= "01110100"; z_correct<="1101010101101000";
        when 8949 => y_in <= "10100010"; x_in <= "01110101"; z_correct<="1101010100001010";
        when 8950 => y_in <= "10100010"; x_in <= "01110110"; z_correct<="1101010010101100";
        when 8951 => y_in <= "10100010"; x_in <= "01110111"; z_correct<="1101010001001110";
        when 8952 => y_in <= "10100010"; x_in <= "01111000"; z_correct<="1101001111110000";
        when 8953 => y_in <= "10100010"; x_in <= "01111001"; z_correct<="1101001110010010";
        when 8954 => y_in <= "10100010"; x_in <= "01111010"; z_correct<="1101001100110100";
        when 8955 => y_in <= "10100010"; x_in <= "01111011"; z_correct<="1101001011010110";
        when 8956 => y_in <= "10100010"; x_in <= "01111100"; z_correct<="1101001001111000";
        when 8957 => y_in <= "10100010"; x_in <= "01111101"; z_correct<="1101001000011010";
        when 8958 => y_in <= "10100010"; x_in <= "01111110"; z_correct<="1101000110111100";
        when 8959 => y_in <= "10100010"; x_in <= "01111111"; z_correct<="1101000101011110";
        when 8960 => y_in <= "10100011"; x_in <= "10000000"; z_correct<="0010111010000000";
        when 8961 => y_in <= "10100011"; x_in <= "10000001"; z_correct<="0010111000100011";
        when 8962 => y_in <= "10100011"; x_in <= "10000010"; z_correct<="0010110111000110";
        when 8963 => y_in <= "10100011"; x_in <= "10000011"; z_correct<="0010110101101001";
        when 8964 => y_in <= "10100011"; x_in <= "10000100"; z_correct<="0010110100001100";
        when 8965 => y_in <= "10100011"; x_in <= "10000101"; z_correct<="0010110010101111";
        when 8966 => y_in <= "10100011"; x_in <= "10000110"; z_correct<="0010110001010010";
        when 8967 => y_in <= "10100011"; x_in <= "10000111"; z_correct<="0010101111110101";
        when 8968 => y_in <= "10100011"; x_in <= "10001000"; z_correct<="0010101110011000";
        when 8969 => y_in <= "10100011"; x_in <= "10001001"; z_correct<="0010101100111011";
        when 8970 => y_in <= "10100011"; x_in <= "10001010"; z_correct<="0010101011011110";
        when 8971 => y_in <= "10100011"; x_in <= "10001011"; z_correct<="0010101010000001";
        when 8972 => y_in <= "10100011"; x_in <= "10001100"; z_correct<="0010101000100100";
        when 8973 => y_in <= "10100011"; x_in <= "10001101"; z_correct<="0010100111000111";
        when 8974 => y_in <= "10100011"; x_in <= "10001110"; z_correct<="0010100101101010";
        when 8975 => y_in <= "10100011"; x_in <= "10001111"; z_correct<="0010100100001101";
        when 8976 => y_in <= "10100011"; x_in <= "10010000"; z_correct<="0010100010110000";
        when 8977 => y_in <= "10100011"; x_in <= "10010001"; z_correct<="0010100001010011";
        when 8978 => y_in <= "10100011"; x_in <= "10010010"; z_correct<="0010011111110110";
        when 8979 => y_in <= "10100011"; x_in <= "10010011"; z_correct<="0010011110011001";
        when 8980 => y_in <= "10100011"; x_in <= "10010100"; z_correct<="0010011100111100";
        when 8981 => y_in <= "10100011"; x_in <= "10010101"; z_correct<="0010011011011111";
        when 8982 => y_in <= "10100011"; x_in <= "10010110"; z_correct<="0010011010000010";
        when 8983 => y_in <= "10100011"; x_in <= "10010111"; z_correct<="0010011000100101";
        when 8984 => y_in <= "10100011"; x_in <= "10011000"; z_correct<="0010010111001000";
        when 8985 => y_in <= "10100011"; x_in <= "10011001"; z_correct<="0010010101101011";
        when 8986 => y_in <= "10100011"; x_in <= "10011010"; z_correct<="0010010100001110";
        when 8987 => y_in <= "10100011"; x_in <= "10011011"; z_correct<="0010010010110001";
        when 8988 => y_in <= "10100011"; x_in <= "10011100"; z_correct<="0010010001010100";
        when 8989 => y_in <= "10100011"; x_in <= "10011101"; z_correct<="0010001111110111";
        when 8990 => y_in <= "10100011"; x_in <= "10011110"; z_correct<="0010001110011010";
        when 8991 => y_in <= "10100011"; x_in <= "10011111"; z_correct<="0010001100111101";
        when 8992 => y_in <= "10100011"; x_in <= "10100000"; z_correct<="0010001011100000";
        when 8993 => y_in <= "10100011"; x_in <= "10100001"; z_correct<="0010001010000011";
        when 8994 => y_in <= "10100011"; x_in <= "10100010"; z_correct<="0010001000100110";
        when 8995 => y_in <= "10100011"; x_in <= "10100011"; z_correct<="0010000111001001";
        when 8996 => y_in <= "10100011"; x_in <= "10100100"; z_correct<="0010000101101100";
        when 8997 => y_in <= "10100011"; x_in <= "10100101"; z_correct<="0010000100001111";
        when 8998 => y_in <= "10100011"; x_in <= "10100110"; z_correct<="0010000010110010";
        when 8999 => y_in <= "10100011"; x_in <= "10100111"; z_correct<="0010000001010101";
        when 9000 => y_in <= "10100011"; x_in <= "10101000"; z_correct<="0001111111111000";
        when 9001 => y_in <= "10100011"; x_in <= "10101001"; z_correct<="0001111110011011";
        when 9002 => y_in <= "10100011"; x_in <= "10101010"; z_correct<="0001111100111110";
        when 9003 => y_in <= "10100011"; x_in <= "10101011"; z_correct<="0001111011100001";
        when 9004 => y_in <= "10100011"; x_in <= "10101100"; z_correct<="0001111010000100";
        when 9005 => y_in <= "10100011"; x_in <= "10101101"; z_correct<="0001111000100111";
        when 9006 => y_in <= "10100011"; x_in <= "10101110"; z_correct<="0001110111001010";
        when 9007 => y_in <= "10100011"; x_in <= "10101111"; z_correct<="0001110101101101";
        when 9008 => y_in <= "10100011"; x_in <= "10110000"; z_correct<="0001110100010000";
        when 9009 => y_in <= "10100011"; x_in <= "10110001"; z_correct<="0001110010110011";
        when 9010 => y_in <= "10100011"; x_in <= "10110010"; z_correct<="0001110001010110";
        when 9011 => y_in <= "10100011"; x_in <= "10110011"; z_correct<="0001101111111001";
        when 9012 => y_in <= "10100011"; x_in <= "10110100"; z_correct<="0001101110011100";
        when 9013 => y_in <= "10100011"; x_in <= "10110101"; z_correct<="0001101100111111";
        when 9014 => y_in <= "10100011"; x_in <= "10110110"; z_correct<="0001101011100010";
        when 9015 => y_in <= "10100011"; x_in <= "10110111"; z_correct<="0001101010000101";
        when 9016 => y_in <= "10100011"; x_in <= "10111000"; z_correct<="0001101000101000";
        when 9017 => y_in <= "10100011"; x_in <= "10111001"; z_correct<="0001100111001011";
        when 9018 => y_in <= "10100011"; x_in <= "10111010"; z_correct<="0001100101101110";
        when 9019 => y_in <= "10100011"; x_in <= "10111011"; z_correct<="0001100100010001";
        when 9020 => y_in <= "10100011"; x_in <= "10111100"; z_correct<="0001100010110100";
        when 9021 => y_in <= "10100011"; x_in <= "10111101"; z_correct<="0001100001010111";
        when 9022 => y_in <= "10100011"; x_in <= "10111110"; z_correct<="0001011111111010";
        when 9023 => y_in <= "10100011"; x_in <= "10111111"; z_correct<="0001011110011101";
        when 9024 => y_in <= "10100011"; x_in <= "11000000"; z_correct<="0001011101000000";
        when 9025 => y_in <= "10100011"; x_in <= "11000001"; z_correct<="0001011011100011";
        when 9026 => y_in <= "10100011"; x_in <= "11000010"; z_correct<="0001011010000110";
        when 9027 => y_in <= "10100011"; x_in <= "11000011"; z_correct<="0001011000101001";
        when 9028 => y_in <= "10100011"; x_in <= "11000100"; z_correct<="0001010111001100";
        when 9029 => y_in <= "10100011"; x_in <= "11000101"; z_correct<="0001010101101111";
        when 9030 => y_in <= "10100011"; x_in <= "11000110"; z_correct<="0001010100010010";
        when 9031 => y_in <= "10100011"; x_in <= "11000111"; z_correct<="0001010010110101";
        when 9032 => y_in <= "10100011"; x_in <= "11001000"; z_correct<="0001010001011000";
        when 9033 => y_in <= "10100011"; x_in <= "11001001"; z_correct<="0001001111111011";
        when 9034 => y_in <= "10100011"; x_in <= "11001010"; z_correct<="0001001110011110";
        when 9035 => y_in <= "10100011"; x_in <= "11001011"; z_correct<="0001001101000001";
        when 9036 => y_in <= "10100011"; x_in <= "11001100"; z_correct<="0001001011100100";
        when 9037 => y_in <= "10100011"; x_in <= "11001101"; z_correct<="0001001010000111";
        when 9038 => y_in <= "10100011"; x_in <= "11001110"; z_correct<="0001001000101010";
        when 9039 => y_in <= "10100011"; x_in <= "11001111"; z_correct<="0001000111001101";
        when 9040 => y_in <= "10100011"; x_in <= "11010000"; z_correct<="0001000101110000";
        when 9041 => y_in <= "10100011"; x_in <= "11010001"; z_correct<="0001000100010011";
        when 9042 => y_in <= "10100011"; x_in <= "11010010"; z_correct<="0001000010110110";
        when 9043 => y_in <= "10100011"; x_in <= "11010011"; z_correct<="0001000001011001";
        when 9044 => y_in <= "10100011"; x_in <= "11010100"; z_correct<="0000111111111100";
        when 9045 => y_in <= "10100011"; x_in <= "11010101"; z_correct<="0000111110011111";
        when 9046 => y_in <= "10100011"; x_in <= "11010110"; z_correct<="0000111101000010";
        when 9047 => y_in <= "10100011"; x_in <= "11010111"; z_correct<="0000111011100101";
        when 9048 => y_in <= "10100011"; x_in <= "11011000"; z_correct<="0000111010001000";
        when 9049 => y_in <= "10100011"; x_in <= "11011001"; z_correct<="0000111000101011";
        when 9050 => y_in <= "10100011"; x_in <= "11011010"; z_correct<="0000110111001110";
        when 9051 => y_in <= "10100011"; x_in <= "11011011"; z_correct<="0000110101110001";
        when 9052 => y_in <= "10100011"; x_in <= "11011100"; z_correct<="0000110100010100";
        when 9053 => y_in <= "10100011"; x_in <= "11011101"; z_correct<="0000110010110111";
        when 9054 => y_in <= "10100011"; x_in <= "11011110"; z_correct<="0000110001011010";
        when 9055 => y_in <= "10100011"; x_in <= "11011111"; z_correct<="0000101111111101";
        when 9056 => y_in <= "10100011"; x_in <= "11100000"; z_correct<="0000101110100000";
        when 9057 => y_in <= "10100011"; x_in <= "11100001"; z_correct<="0000101101000011";
        when 9058 => y_in <= "10100011"; x_in <= "11100010"; z_correct<="0000101011100110";
        when 9059 => y_in <= "10100011"; x_in <= "11100011"; z_correct<="0000101010001001";
        when 9060 => y_in <= "10100011"; x_in <= "11100100"; z_correct<="0000101000101100";
        when 9061 => y_in <= "10100011"; x_in <= "11100101"; z_correct<="0000100111001111";
        when 9062 => y_in <= "10100011"; x_in <= "11100110"; z_correct<="0000100101110010";
        when 9063 => y_in <= "10100011"; x_in <= "11100111"; z_correct<="0000100100010101";
        when 9064 => y_in <= "10100011"; x_in <= "11101000"; z_correct<="0000100010111000";
        when 9065 => y_in <= "10100011"; x_in <= "11101001"; z_correct<="0000100001011011";
        when 9066 => y_in <= "10100011"; x_in <= "11101010"; z_correct<="0000011111111110";
        when 9067 => y_in <= "10100011"; x_in <= "11101011"; z_correct<="0000011110100001";
        when 9068 => y_in <= "10100011"; x_in <= "11101100"; z_correct<="0000011101000100";
        when 9069 => y_in <= "10100011"; x_in <= "11101101"; z_correct<="0000011011100111";
        when 9070 => y_in <= "10100011"; x_in <= "11101110"; z_correct<="0000011010001010";
        when 9071 => y_in <= "10100011"; x_in <= "11101111"; z_correct<="0000011000101101";
        when 9072 => y_in <= "10100011"; x_in <= "11110000"; z_correct<="0000010111010000";
        when 9073 => y_in <= "10100011"; x_in <= "11110001"; z_correct<="0000010101110011";
        when 9074 => y_in <= "10100011"; x_in <= "11110010"; z_correct<="0000010100010110";
        when 9075 => y_in <= "10100011"; x_in <= "11110011"; z_correct<="0000010010111001";
        when 9076 => y_in <= "10100011"; x_in <= "11110100"; z_correct<="0000010001011100";
        when 9077 => y_in <= "10100011"; x_in <= "11110101"; z_correct<="0000001111111111";
        when 9078 => y_in <= "10100011"; x_in <= "11110110"; z_correct<="0000001110100010";
        when 9079 => y_in <= "10100011"; x_in <= "11110111"; z_correct<="0000001101000101";
        when 9080 => y_in <= "10100011"; x_in <= "11111000"; z_correct<="0000001011101000";
        when 9081 => y_in <= "10100011"; x_in <= "11111001"; z_correct<="0000001010001011";
        when 9082 => y_in <= "10100011"; x_in <= "11111010"; z_correct<="0000001000101110";
        when 9083 => y_in <= "10100011"; x_in <= "11111011"; z_correct<="0000000111010001";
        when 9084 => y_in <= "10100011"; x_in <= "11111100"; z_correct<="0000000101110100";
        when 9085 => y_in <= "10100011"; x_in <= "11111101"; z_correct<="0000000100010111";
        when 9086 => y_in <= "10100011"; x_in <= "11111110"; z_correct<="0000000010111010";
        when 9087 => y_in <= "10100011"; x_in <= "11111111"; z_correct<="0000000001011101";
        when 9088 => y_in <= "10100011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 9089 => y_in <= "10100011"; x_in <= "00000001"; z_correct<="1111111110100011";
        when 9090 => y_in <= "10100011"; x_in <= "00000010"; z_correct<="1111111101000110";
        when 9091 => y_in <= "10100011"; x_in <= "00000011"; z_correct<="1111111011101001";
        when 9092 => y_in <= "10100011"; x_in <= "00000100"; z_correct<="1111111010001100";
        when 9093 => y_in <= "10100011"; x_in <= "00000101"; z_correct<="1111111000101111";
        when 9094 => y_in <= "10100011"; x_in <= "00000110"; z_correct<="1111110111010010";
        when 9095 => y_in <= "10100011"; x_in <= "00000111"; z_correct<="1111110101110101";
        when 9096 => y_in <= "10100011"; x_in <= "00001000"; z_correct<="1111110100011000";
        when 9097 => y_in <= "10100011"; x_in <= "00001001"; z_correct<="1111110010111011";
        when 9098 => y_in <= "10100011"; x_in <= "00001010"; z_correct<="1111110001011110";
        when 9099 => y_in <= "10100011"; x_in <= "00001011"; z_correct<="1111110000000001";
        when 9100 => y_in <= "10100011"; x_in <= "00001100"; z_correct<="1111101110100100";
        when 9101 => y_in <= "10100011"; x_in <= "00001101"; z_correct<="1111101101000111";
        when 9102 => y_in <= "10100011"; x_in <= "00001110"; z_correct<="1111101011101010";
        when 9103 => y_in <= "10100011"; x_in <= "00001111"; z_correct<="1111101010001101";
        when 9104 => y_in <= "10100011"; x_in <= "00010000"; z_correct<="1111101000110000";
        when 9105 => y_in <= "10100011"; x_in <= "00010001"; z_correct<="1111100111010011";
        when 9106 => y_in <= "10100011"; x_in <= "00010010"; z_correct<="1111100101110110";
        when 9107 => y_in <= "10100011"; x_in <= "00010011"; z_correct<="1111100100011001";
        when 9108 => y_in <= "10100011"; x_in <= "00010100"; z_correct<="1111100010111100";
        when 9109 => y_in <= "10100011"; x_in <= "00010101"; z_correct<="1111100001011111";
        when 9110 => y_in <= "10100011"; x_in <= "00010110"; z_correct<="1111100000000010";
        when 9111 => y_in <= "10100011"; x_in <= "00010111"; z_correct<="1111011110100101";
        when 9112 => y_in <= "10100011"; x_in <= "00011000"; z_correct<="1111011101001000";
        when 9113 => y_in <= "10100011"; x_in <= "00011001"; z_correct<="1111011011101011";
        when 9114 => y_in <= "10100011"; x_in <= "00011010"; z_correct<="1111011010001110";
        when 9115 => y_in <= "10100011"; x_in <= "00011011"; z_correct<="1111011000110001";
        when 9116 => y_in <= "10100011"; x_in <= "00011100"; z_correct<="1111010111010100";
        when 9117 => y_in <= "10100011"; x_in <= "00011101"; z_correct<="1111010101110111";
        when 9118 => y_in <= "10100011"; x_in <= "00011110"; z_correct<="1111010100011010";
        when 9119 => y_in <= "10100011"; x_in <= "00011111"; z_correct<="1111010010111101";
        when 9120 => y_in <= "10100011"; x_in <= "00100000"; z_correct<="1111010001100000";
        when 9121 => y_in <= "10100011"; x_in <= "00100001"; z_correct<="1111010000000011";
        when 9122 => y_in <= "10100011"; x_in <= "00100010"; z_correct<="1111001110100110";
        when 9123 => y_in <= "10100011"; x_in <= "00100011"; z_correct<="1111001101001001";
        when 9124 => y_in <= "10100011"; x_in <= "00100100"; z_correct<="1111001011101100";
        when 9125 => y_in <= "10100011"; x_in <= "00100101"; z_correct<="1111001010001111";
        when 9126 => y_in <= "10100011"; x_in <= "00100110"; z_correct<="1111001000110010";
        when 9127 => y_in <= "10100011"; x_in <= "00100111"; z_correct<="1111000111010101";
        when 9128 => y_in <= "10100011"; x_in <= "00101000"; z_correct<="1111000101111000";
        when 9129 => y_in <= "10100011"; x_in <= "00101001"; z_correct<="1111000100011011";
        when 9130 => y_in <= "10100011"; x_in <= "00101010"; z_correct<="1111000010111110";
        when 9131 => y_in <= "10100011"; x_in <= "00101011"; z_correct<="1111000001100001";
        when 9132 => y_in <= "10100011"; x_in <= "00101100"; z_correct<="1111000000000100";
        when 9133 => y_in <= "10100011"; x_in <= "00101101"; z_correct<="1110111110100111";
        when 9134 => y_in <= "10100011"; x_in <= "00101110"; z_correct<="1110111101001010";
        when 9135 => y_in <= "10100011"; x_in <= "00101111"; z_correct<="1110111011101101";
        when 9136 => y_in <= "10100011"; x_in <= "00110000"; z_correct<="1110111010010000";
        when 9137 => y_in <= "10100011"; x_in <= "00110001"; z_correct<="1110111000110011";
        when 9138 => y_in <= "10100011"; x_in <= "00110010"; z_correct<="1110110111010110";
        when 9139 => y_in <= "10100011"; x_in <= "00110011"; z_correct<="1110110101111001";
        when 9140 => y_in <= "10100011"; x_in <= "00110100"; z_correct<="1110110100011100";
        when 9141 => y_in <= "10100011"; x_in <= "00110101"; z_correct<="1110110010111111";
        when 9142 => y_in <= "10100011"; x_in <= "00110110"; z_correct<="1110110001100010";
        when 9143 => y_in <= "10100011"; x_in <= "00110111"; z_correct<="1110110000000101";
        when 9144 => y_in <= "10100011"; x_in <= "00111000"; z_correct<="1110101110101000";
        when 9145 => y_in <= "10100011"; x_in <= "00111001"; z_correct<="1110101101001011";
        when 9146 => y_in <= "10100011"; x_in <= "00111010"; z_correct<="1110101011101110";
        when 9147 => y_in <= "10100011"; x_in <= "00111011"; z_correct<="1110101010010001";
        when 9148 => y_in <= "10100011"; x_in <= "00111100"; z_correct<="1110101000110100";
        when 9149 => y_in <= "10100011"; x_in <= "00111101"; z_correct<="1110100111010111";
        when 9150 => y_in <= "10100011"; x_in <= "00111110"; z_correct<="1110100101111010";
        when 9151 => y_in <= "10100011"; x_in <= "00111111"; z_correct<="1110100100011101";
        when 9152 => y_in <= "10100011"; x_in <= "01000000"; z_correct<="1110100011000000";
        when 9153 => y_in <= "10100011"; x_in <= "01000001"; z_correct<="1110100001100011";
        when 9154 => y_in <= "10100011"; x_in <= "01000010"; z_correct<="1110100000000110";
        when 9155 => y_in <= "10100011"; x_in <= "01000011"; z_correct<="1110011110101001";
        when 9156 => y_in <= "10100011"; x_in <= "01000100"; z_correct<="1110011101001100";
        when 9157 => y_in <= "10100011"; x_in <= "01000101"; z_correct<="1110011011101111";
        when 9158 => y_in <= "10100011"; x_in <= "01000110"; z_correct<="1110011010010010";
        when 9159 => y_in <= "10100011"; x_in <= "01000111"; z_correct<="1110011000110101";
        when 9160 => y_in <= "10100011"; x_in <= "01001000"; z_correct<="1110010111011000";
        when 9161 => y_in <= "10100011"; x_in <= "01001001"; z_correct<="1110010101111011";
        when 9162 => y_in <= "10100011"; x_in <= "01001010"; z_correct<="1110010100011110";
        when 9163 => y_in <= "10100011"; x_in <= "01001011"; z_correct<="1110010011000001";
        when 9164 => y_in <= "10100011"; x_in <= "01001100"; z_correct<="1110010001100100";
        when 9165 => y_in <= "10100011"; x_in <= "01001101"; z_correct<="1110010000000111";
        when 9166 => y_in <= "10100011"; x_in <= "01001110"; z_correct<="1110001110101010";
        when 9167 => y_in <= "10100011"; x_in <= "01001111"; z_correct<="1110001101001101";
        when 9168 => y_in <= "10100011"; x_in <= "01010000"; z_correct<="1110001011110000";
        when 9169 => y_in <= "10100011"; x_in <= "01010001"; z_correct<="1110001010010011";
        when 9170 => y_in <= "10100011"; x_in <= "01010010"; z_correct<="1110001000110110";
        when 9171 => y_in <= "10100011"; x_in <= "01010011"; z_correct<="1110000111011001";
        when 9172 => y_in <= "10100011"; x_in <= "01010100"; z_correct<="1110000101111100";
        when 9173 => y_in <= "10100011"; x_in <= "01010101"; z_correct<="1110000100011111";
        when 9174 => y_in <= "10100011"; x_in <= "01010110"; z_correct<="1110000011000010";
        when 9175 => y_in <= "10100011"; x_in <= "01010111"; z_correct<="1110000001100101";
        when 9176 => y_in <= "10100011"; x_in <= "01011000"; z_correct<="1110000000001000";
        when 9177 => y_in <= "10100011"; x_in <= "01011001"; z_correct<="1101111110101011";
        when 9178 => y_in <= "10100011"; x_in <= "01011010"; z_correct<="1101111101001110";
        when 9179 => y_in <= "10100011"; x_in <= "01011011"; z_correct<="1101111011110001";
        when 9180 => y_in <= "10100011"; x_in <= "01011100"; z_correct<="1101111010010100";
        when 9181 => y_in <= "10100011"; x_in <= "01011101"; z_correct<="1101111000110111";
        when 9182 => y_in <= "10100011"; x_in <= "01011110"; z_correct<="1101110111011010";
        when 9183 => y_in <= "10100011"; x_in <= "01011111"; z_correct<="1101110101111101";
        when 9184 => y_in <= "10100011"; x_in <= "01100000"; z_correct<="1101110100100000";
        when 9185 => y_in <= "10100011"; x_in <= "01100001"; z_correct<="1101110011000011";
        when 9186 => y_in <= "10100011"; x_in <= "01100010"; z_correct<="1101110001100110";
        when 9187 => y_in <= "10100011"; x_in <= "01100011"; z_correct<="1101110000001001";
        when 9188 => y_in <= "10100011"; x_in <= "01100100"; z_correct<="1101101110101100";
        when 9189 => y_in <= "10100011"; x_in <= "01100101"; z_correct<="1101101101001111";
        when 9190 => y_in <= "10100011"; x_in <= "01100110"; z_correct<="1101101011110010";
        when 9191 => y_in <= "10100011"; x_in <= "01100111"; z_correct<="1101101010010101";
        when 9192 => y_in <= "10100011"; x_in <= "01101000"; z_correct<="1101101000111000";
        when 9193 => y_in <= "10100011"; x_in <= "01101001"; z_correct<="1101100111011011";
        when 9194 => y_in <= "10100011"; x_in <= "01101010"; z_correct<="1101100101111110";
        when 9195 => y_in <= "10100011"; x_in <= "01101011"; z_correct<="1101100100100001";
        when 9196 => y_in <= "10100011"; x_in <= "01101100"; z_correct<="1101100011000100";
        when 9197 => y_in <= "10100011"; x_in <= "01101101"; z_correct<="1101100001100111";
        when 9198 => y_in <= "10100011"; x_in <= "01101110"; z_correct<="1101100000001010";
        when 9199 => y_in <= "10100011"; x_in <= "01101111"; z_correct<="1101011110101101";
        when 9200 => y_in <= "10100011"; x_in <= "01110000"; z_correct<="1101011101010000";
        when 9201 => y_in <= "10100011"; x_in <= "01110001"; z_correct<="1101011011110011";
        when 9202 => y_in <= "10100011"; x_in <= "01110010"; z_correct<="1101011010010110";
        when 9203 => y_in <= "10100011"; x_in <= "01110011"; z_correct<="1101011000111001";
        when 9204 => y_in <= "10100011"; x_in <= "01110100"; z_correct<="1101010111011100";
        when 9205 => y_in <= "10100011"; x_in <= "01110101"; z_correct<="1101010101111111";
        when 9206 => y_in <= "10100011"; x_in <= "01110110"; z_correct<="1101010100100010";
        when 9207 => y_in <= "10100011"; x_in <= "01110111"; z_correct<="1101010011000101";
        when 9208 => y_in <= "10100011"; x_in <= "01111000"; z_correct<="1101010001101000";
        when 9209 => y_in <= "10100011"; x_in <= "01111001"; z_correct<="1101010000001011";
        when 9210 => y_in <= "10100011"; x_in <= "01111010"; z_correct<="1101001110101110";
        when 9211 => y_in <= "10100011"; x_in <= "01111011"; z_correct<="1101001101010001";
        when 9212 => y_in <= "10100011"; x_in <= "01111100"; z_correct<="1101001011110100";
        when 9213 => y_in <= "10100011"; x_in <= "01111101"; z_correct<="1101001010010111";
        when 9214 => y_in <= "10100011"; x_in <= "01111110"; z_correct<="1101001000111010";
        when 9215 => y_in <= "10100011"; x_in <= "01111111"; z_correct<="1101000111011101";
        when 9216 => y_in <= "10100100"; x_in <= "10000000"; z_correct<="0010111000000000";
        when 9217 => y_in <= "10100100"; x_in <= "10000001"; z_correct<="0010110110100100";
        when 9218 => y_in <= "10100100"; x_in <= "10000010"; z_correct<="0010110101001000";
        when 9219 => y_in <= "10100100"; x_in <= "10000011"; z_correct<="0010110011101100";
        when 9220 => y_in <= "10100100"; x_in <= "10000100"; z_correct<="0010110010010000";
        when 9221 => y_in <= "10100100"; x_in <= "10000101"; z_correct<="0010110000110100";
        when 9222 => y_in <= "10100100"; x_in <= "10000110"; z_correct<="0010101111011000";
        when 9223 => y_in <= "10100100"; x_in <= "10000111"; z_correct<="0010101101111100";
        when 9224 => y_in <= "10100100"; x_in <= "10001000"; z_correct<="0010101100100000";
        when 9225 => y_in <= "10100100"; x_in <= "10001001"; z_correct<="0010101011000100";
        when 9226 => y_in <= "10100100"; x_in <= "10001010"; z_correct<="0010101001101000";
        when 9227 => y_in <= "10100100"; x_in <= "10001011"; z_correct<="0010101000001100";
        when 9228 => y_in <= "10100100"; x_in <= "10001100"; z_correct<="0010100110110000";
        when 9229 => y_in <= "10100100"; x_in <= "10001101"; z_correct<="0010100101010100";
        when 9230 => y_in <= "10100100"; x_in <= "10001110"; z_correct<="0010100011111000";
        when 9231 => y_in <= "10100100"; x_in <= "10001111"; z_correct<="0010100010011100";
        when 9232 => y_in <= "10100100"; x_in <= "10010000"; z_correct<="0010100001000000";
        when 9233 => y_in <= "10100100"; x_in <= "10010001"; z_correct<="0010011111100100";
        when 9234 => y_in <= "10100100"; x_in <= "10010010"; z_correct<="0010011110001000";
        when 9235 => y_in <= "10100100"; x_in <= "10010011"; z_correct<="0010011100101100";
        when 9236 => y_in <= "10100100"; x_in <= "10010100"; z_correct<="0010011011010000";
        when 9237 => y_in <= "10100100"; x_in <= "10010101"; z_correct<="0010011001110100";
        when 9238 => y_in <= "10100100"; x_in <= "10010110"; z_correct<="0010011000011000";
        when 9239 => y_in <= "10100100"; x_in <= "10010111"; z_correct<="0010010110111100";
        when 9240 => y_in <= "10100100"; x_in <= "10011000"; z_correct<="0010010101100000";
        when 9241 => y_in <= "10100100"; x_in <= "10011001"; z_correct<="0010010100000100";
        when 9242 => y_in <= "10100100"; x_in <= "10011010"; z_correct<="0010010010101000";
        when 9243 => y_in <= "10100100"; x_in <= "10011011"; z_correct<="0010010001001100";
        when 9244 => y_in <= "10100100"; x_in <= "10011100"; z_correct<="0010001111110000";
        when 9245 => y_in <= "10100100"; x_in <= "10011101"; z_correct<="0010001110010100";
        when 9246 => y_in <= "10100100"; x_in <= "10011110"; z_correct<="0010001100111000";
        when 9247 => y_in <= "10100100"; x_in <= "10011111"; z_correct<="0010001011011100";
        when 9248 => y_in <= "10100100"; x_in <= "10100000"; z_correct<="0010001010000000";
        when 9249 => y_in <= "10100100"; x_in <= "10100001"; z_correct<="0010001000100100";
        when 9250 => y_in <= "10100100"; x_in <= "10100010"; z_correct<="0010000111001000";
        when 9251 => y_in <= "10100100"; x_in <= "10100011"; z_correct<="0010000101101100";
        when 9252 => y_in <= "10100100"; x_in <= "10100100"; z_correct<="0010000100010000";
        when 9253 => y_in <= "10100100"; x_in <= "10100101"; z_correct<="0010000010110100";
        when 9254 => y_in <= "10100100"; x_in <= "10100110"; z_correct<="0010000001011000";
        when 9255 => y_in <= "10100100"; x_in <= "10100111"; z_correct<="0001111111111100";
        when 9256 => y_in <= "10100100"; x_in <= "10101000"; z_correct<="0001111110100000";
        when 9257 => y_in <= "10100100"; x_in <= "10101001"; z_correct<="0001111101000100";
        when 9258 => y_in <= "10100100"; x_in <= "10101010"; z_correct<="0001111011101000";
        when 9259 => y_in <= "10100100"; x_in <= "10101011"; z_correct<="0001111010001100";
        when 9260 => y_in <= "10100100"; x_in <= "10101100"; z_correct<="0001111000110000";
        when 9261 => y_in <= "10100100"; x_in <= "10101101"; z_correct<="0001110111010100";
        when 9262 => y_in <= "10100100"; x_in <= "10101110"; z_correct<="0001110101111000";
        when 9263 => y_in <= "10100100"; x_in <= "10101111"; z_correct<="0001110100011100";
        when 9264 => y_in <= "10100100"; x_in <= "10110000"; z_correct<="0001110011000000";
        when 9265 => y_in <= "10100100"; x_in <= "10110001"; z_correct<="0001110001100100";
        when 9266 => y_in <= "10100100"; x_in <= "10110010"; z_correct<="0001110000001000";
        when 9267 => y_in <= "10100100"; x_in <= "10110011"; z_correct<="0001101110101100";
        when 9268 => y_in <= "10100100"; x_in <= "10110100"; z_correct<="0001101101010000";
        when 9269 => y_in <= "10100100"; x_in <= "10110101"; z_correct<="0001101011110100";
        when 9270 => y_in <= "10100100"; x_in <= "10110110"; z_correct<="0001101010011000";
        when 9271 => y_in <= "10100100"; x_in <= "10110111"; z_correct<="0001101000111100";
        when 9272 => y_in <= "10100100"; x_in <= "10111000"; z_correct<="0001100111100000";
        when 9273 => y_in <= "10100100"; x_in <= "10111001"; z_correct<="0001100110000100";
        when 9274 => y_in <= "10100100"; x_in <= "10111010"; z_correct<="0001100100101000";
        when 9275 => y_in <= "10100100"; x_in <= "10111011"; z_correct<="0001100011001100";
        when 9276 => y_in <= "10100100"; x_in <= "10111100"; z_correct<="0001100001110000";
        when 9277 => y_in <= "10100100"; x_in <= "10111101"; z_correct<="0001100000010100";
        when 9278 => y_in <= "10100100"; x_in <= "10111110"; z_correct<="0001011110111000";
        when 9279 => y_in <= "10100100"; x_in <= "10111111"; z_correct<="0001011101011100";
        when 9280 => y_in <= "10100100"; x_in <= "11000000"; z_correct<="0001011100000000";
        when 9281 => y_in <= "10100100"; x_in <= "11000001"; z_correct<="0001011010100100";
        when 9282 => y_in <= "10100100"; x_in <= "11000010"; z_correct<="0001011001001000";
        when 9283 => y_in <= "10100100"; x_in <= "11000011"; z_correct<="0001010111101100";
        when 9284 => y_in <= "10100100"; x_in <= "11000100"; z_correct<="0001010110010000";
        when 9285 => y_in <= "10100100"; x_in <= "11000101"; z_correct<="0001010100110100";
        when 9286 => y_in <= "10100100"; x_in <= "11000110"; z_correct<="0001010011011000";
        when 9287 => y_in <= "10100100"; x_in <= "11000111"; z_correct<="0001010001111100";
        when 9288 => y_in <= "10100100"; x_in <= "11001000"; z_correct<="0001010000100000";
        when 9289 => y_in <= "10100100"; x_in <= "11001001"; z_correct<="0001001111000100";
        when 9290 => y_in <= "10100100"; x_in <= "11001010"; z_correct<="0001001101101000";
        when 9291 => y_in <= "10100100"; x_in <= "11001011"; z_correct<="0001001100001100";
        when 9292 => y_in <= "10100100"; x_in <= "11001100"; z_correct<="0001001010110000";
        when 9293 => y_in <= "10100100"; x_in <= "11001101"; z_correct<="0001001001010100";
        when 9294 => y_in <= "10100100"; x_in <= "11001110"; z_correct<="0001000111111000";
        when 9295 => y_in <= "10100100"; x_in <= "11001111"; z_correct<="0001000110011100";
        when 9296 => y_in <= "10100100"; x_in <= "11010000"; z_correct<="0001000101000000";
        when 9297 => y_in <= "10100100"; x_in <= "11010001"; z_correct<="0001000011100100";
        when 9298 => y_in <= "10100100"; x_in <= "11010010"; z_correct<="0001000010001000";
        when 9299 => y_in <= "10100100"; x_in <= "11010011"; z_correct<="0001000000101100";
        when 9300 => y_in <= "10100100"; x_in <= "11010100"; z_correct<="0000111111010000";
        when 9301 => y_in <= "10100100"; x_in <= "11010101"; z_correct<="0000111101110100";
        when 9302 => y_in <= "10100100"; x_in <= "11010110"; z_correct<="0000111100011000";
        when 9303 => y_in <= "10100100"; x_in <= "11010111"; z_correct<="0000111010111100";
        when 9304 => y_in <= "10100100"; x_in <= "11011000"; z_correct<="0000111001100000";
        when 9305 => y_in <= "10100100"; x_in <= "11011001"; z_correct<="0000111000000100";
        when 9306 => y_in <= "10100100"; x_in <= "11011010"; z_correct<="0000110110101000";
        when 9307 => y_in <= "10100100"; x_in <= "11011011"; z_correct<="0000110101001100";
        when 9308 => y_in <= "10100100"; x_in <= "11011100"; z_correct<="0000110011110000";
        when 9309 => y_in <= "10100100"; x_in <= "11011101"; z_correct<="0000110010010100";
        when 9310 => y_in <= "10100100"; x_in <= "11011110"; z_correct<="0000110000111000";
        when 9311 => y_in <= "10100100"; x_in <= "11011111"; z_correct<="0000101111011100";
        when 9312 => y_in <= "10100100"; x_in <= "11100000"; z_correct<="0000101110000000";
        when 9313 => y_in <= "10100100"; x_in <= "11100001"; z_correct<="0000101100100100";
        when 9314 => y_in <= "10100100"; x_in <= "11100010"; z_correct<="0000101011001000";
        when 9315 => y_in <= "10100100"; x_in <= "11100011"; z_correct<="0000101001101100";
        when 9316 => y_in <= "10100100"; x_in <= "11100100"; z_correct<="0000101000010000";
        when 9317 => y_in <= "10100100"; x_in <= "11100101"; z_correct<="0000100110110100";
        when 9318 => y_in <= "10100100"; x_in <= "11100110"; z_correct<="0000100101011000";
        when 9319 => y_in <= "10100100"; x_in <= "11100111"; z_correct<="0000100011111100";
        when 9320 => y_in <= "10100100"; x_in <= "11101000"; z_correct<="0000100010100000";
        when 9321 => y_in <= "10100100"; x_in <= "11101001"; z_correct<="0000100001000100";
        when 9322 => y_in <= "10100100"; x_in <= "11101010"; z_correct<="0000011111101000";
        when 9323 => y_in <= "10100100"; x_in <= "11101011"; z_correct<="0000011110001100";
        when 9324 => y_in <= "10100100"; x_in <= "11101100"; z_correct<="0000011100110000";
        when 9325 => y_in <= "10100100"; x_in <= "11101101"; z_correct<="0000011011010100";
        when 9326 => y_in <= "10100100"; x_in <= "11101110"; z_correct<="0000011001111000";
        when 9327 => y_in <= "10100100"; x_in <= "11101111"; z_correct<="0000011000011100";
        when 9328 => y_in <= "10100100"; x_in <= "11110000"; z_correct<="0000010111000000";
        when 9329 => y_in <= "10100100"; x_in <= "11110001"; z_correct<="0000010101100100";
        when 9330 => y_in <= "10100100"; x_in <= "11110010"; z_correct<="0000010100001000";
        when 9331 => y_in <= "10100100"; x_in <= "11110011"; z_correct<="0000010010101100";
        when 9332 => y_in <= "10100100"; x_in <= "11110100"; z_correct<="0000010001010000";
        when 9333 => y_in <= "10100100"; x_in <= "11110101"; z_correct<="0000001111110100";
        when 9334 => y_in <= "10100100"; x_in <= "11110110"; z_correct<="0000001110011000";
        when 9335 => y_in <= "10100100"; x_in <= "11110111"; z_correct<="0000001100111100";
        when 9336 => y_in <= "10100100"; x_in <= "11111000"; z_correct<="0000001011100000";
        when 9337 => y_in <= "10100100"; x_in <= "11111001"; z_correct<="0000001010000100";
        when 9338 => y_in <= "10100100"; x_in <= "11111010"; z_correct<="0000001000101000";
        when 9339 => y_in <= "10100100"; x_in <= "11111011"; z_correct<="0000000111001100";
        when 9340 => y_in <= "10100100"; x_in <= "11111100"; z_correct<="0000000101110000";
        when 9341 => y_in <= "10100100"; x_in <= "11111101"; z_correct<="0000000100010100";
        when 9342 => y_in <= "10100100"; x_in <= "11111110"; z_correct<="0000000010111000";
        when 9343 => y_in <= "10100100"; x_in <= "11111111"; z_correct<="0000000001011100";
        when 9344 => y_in <= "10100100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 9345 => y_in <= "10100100"; x_in <= "00000001"; z_correct<="1111111110100100";
        when 9346 => y_in <= "10100100"; x_in <= "00000010"; z_correct<="1111111101001000";
        when 9347 => y_in <= "10100100"; x_in <= "00000011"; z_correct<="1111111011101100";
        when 9348 => y_in <= "10100100"; x_in <= "00000100"; z_correct<="1111111010010000";
        when 9349 => y_in <= "10100100"; x_in <= "00000101"; z_correct<="1111111000110100";
        when 9350 => y_in <= "10100100"; x_in <= "00000110"; z_correct<="1111110111011000";
        when 9351 => y_in <= "10100100"; x_in <= "00000111"; z_correct<="1111110101111100";
        when 9352 => y_in <= "10100100"; x_in <= "00001000"; z_correct<="1111110100100000";
        when 9353 => y_in <= "10100100"; x_in <= "00001001"; z_correct<="1111110011000100";
        when 9354 => y_in <= "10100100"; x_in <= "00001010"; z_correct<="1111110001101000";
        when 9355 => y_in <= "10100100"; x_in <= "00001011"; z_correct<="1111110000001100";
        when 9356 => y_in <= "10100100"; x_in <= "00001100"; z_correct<="1111101110110000";
        when 9357 => y_in <= "10100100"; x_in <= "00001101"; z_correct<="1111101101010100";
        when 9358 => y_in <= "10100100"; x_in <= "00001110"; z_correct<="1111101011111000";
        when 9359 => y_in <= "10100100"; x_in <= "00001111"; z_correct<="1111101010011100";
        when 9360 => y_in <= "10100100"; x_in <= "00010000"; z_correct<="1111101001000000";
        when 9361 => y_in <= "10100100"; x_in <= "00010001"; z_correct<="1111100111100100";
        when 9362 => y_in <= "10100100"; x_in <= "00010010"; z_correct<="1111100110001000";
        when 9363 => y_in <= "10100100"; x_in <= "00010011"; z_correct<="1111100100101100";
        when 9364 => y_in <= "10100100"; x_in <= "00010100"; z_correct<="1111100011010000";
        when 9365 => y_in <= "10100100"; x_in <= "00010101"; z_correct<="1111100001110100";
        when 9366 => y_in <= "10100100"; x_in <= "00010110"; z_correct<="1111100000011000";
        when 9367 => y_in <= "10100100"; x_in <= "00010111"; z_correct<="1111011110111100";
        when 9368 => y_in <= "10100100"; x_in <= "00011000"; z_correct<="1111011101100000";
        when 9369 => y_in <= "10100100"; x_in <= "00011001"; z_correct<="1111011100000100";
        when 9370 => y_in <= "10100100"; x_in <= "00011010"; z_correct<="1111011010101000";
        when 9371 => y_in <= "10100100"; x_in <= "00011011"; z_correct<="1111011001001100";
        when 9372 => y_in <= "10100100"; x_in <= "00011100"; z_correct<="1111010111110000";
        when 9373 => y_in <= "10100100"; x_in <= "00011101"; z_correct<="1111010110010100";
        when 9374 => y_in <= "10100100"; x_in <= "00011110"; z_correct<="1111010100111000";
        when 9375 => y_in <= "10100100"; x_in <= "00011111"; z_correct<="1111010011011100";
        when 9376 => y_in <= "10100100"; x_in <= "00100000"; z_correct<="1111010010000000";
        when 9377 => y_in <= "10100100"; x_in <= "00100001"; z_correct<="1111010000100100";
        when 9378 => y_in <= "10100100"; x_in <= "00100010"; z_correct<="1111001111001000";
        when 9379 => y_in <= "10100100"; x_in <= "00100011"; z_correct<="1111001101101100";
        when 9380 => y_in <= "10100100"; x_in <= "00100100"; z_correct<="1111001100010000";
        when 9381 => y_in <= "10100100"; x_in <= "00100101"; z_correct<="1111001010110100";
        when 9382 => y_in <= "10100100"; x_in <= "00100110"; z_correct<="1111001001011000";
        when 9383 => y_in <= "10100100"; x_in <= "00100111"; z_correct<="1111000111111100";
        when 9384 => y_in <= "10100100"; x_in <= "00101000"; z_correct<="1111000110100000";
        when 9385 => y_in <= "10100100"; x_in <= "00101001"; z_correct<="1111000101000100";
        when 9386 => y_in <= "10100100"; x_in <= "00101010"; z_correct<="1111000011101000";
        when 9387 => y_in <= "10100100"; x_in <= "00101011"; z_correct<="1111000010001100";
        when 9388 => y_in <= "10100100"; x_in <= "00101100"; z_correct<="1111000000110000";
        when 9389 => y_in <= "10100100"; x_in <= "00101101"; z_correct<="1110111111010100";
        when 9390 => y_in <= "10100100"; x_in <= "00101110"; z_correct<="1110111101111000";
        when 9391 => y_in <= "10100100"; x_in <= "00101111"; z_correct<="1110111100011100";
        when 9392 => y_in <= "10100100"; x_in <= "00110000"; z_correct<="1110111011000000";
        when 9393 => y_in <= "10100100"; x_in <= "00110001"; z_correct<="1110111001100100";
        when 9394 => y_in <= "10100100"; x_in <= "00110010"; z_correct<="1110111000001000";
        when 9395 => y_in <= "10100100"; x_in <= "00110011"; z_correct<="1110110110101100";
        when 9396 => y_in <= "10100100"; x_in <= "00110100"; z_correct<="1110110101010000";
        when 9397 => y_in <= "10100100"; x_in <= "00110101"; z_correct<="1110110011110100";
        when 9398 => y_in <= "10100100"; x_in <= "00110110"; z_correct<="1110110010011000";
        when 9399 => y_in <= "10100100"; x_in <= "00110111"; z_correct<="1110110000111100";
        when 9400 => y_in <= "10100100"; x_in <= "00111000"; z_correct<="1110101111100000";
        when 9401 => y_in <= "10100100"; x_in <= "00111001"; z_correct<="1110101110000100";
        when 9402 => y_in <= "10100100"; x_in <= "00111010"; z_correct<="1110101100101000";
        when 9403 => y_in <= "10100100"; x_in <= "00111011"; z_correct<="1110101011001100";
        when 9404 => y_in <= "10100100"; x_in <= "00111100"; z_correct<="1110101001110000";
        when 9405 => y_in <= "10100100"; x_in <= "00111101"; z_correct<="1110101000010100";
        when 9406 => y_in <= "10100100"; x_in <= "00111110"; z_correct<="1110100110111000";
        when 9407 => y_in <= "10100100"; x_in <= "00111111"; z_correct<="1110100101011100";
        when 9408 => y_in <= "10100100"; x_in <= "01000000"; z_correct<="1110100100000000";
        when 9409 => y_in <= "10100100"; x_in <= "01000001"; z_correct<="1110100010100100";
        when 9410 => y_in <= "10100100"; x_in <= "01000010"; z_correct<="1110100001001000";
        when 9411 => y_in <= "10100100"; x_in <= "01000011"; z_correct<="1110011111101100";
        when 9412 => y_in <= "10100100"; x_in <= "01000100"; z_correct<="1110011110010000";
        when 9413 => y_in <= "10100100"; x_in <= "01000101"; z_correct<="1110011100110100";
        when 9414 => y_in <= "10100100"; x_in <= "01000110"; z_correct<="1110011011011000";
        when 9415 => y_in <= "10100100"; x_in <= "01000111"; z_correct<="1110011001111100";
        when 9416 => y_in <= "10100100"; x_in <= "01001000"; z_correct<="1110011000100000";
        when 9417 => y_in <= "10100100"; x_in <= "01001001"; z_correct<="1110010111000100";
        when 9418 => y_in <= "10100100"; x_in <= "01001010"; z_correct<="1110010101101000";
        when 9419 => y_in <= "10100100"; x_in <= "01001011"; z_correct<="1110010100001100";
        when 9420 => y_in <= "10100100"; x_in <= "01001100"; z_correct<="1110010010110000";
        when 9421 => y_in <= "10100100"; x_in <= "01001101"; z_correct<="1110010001010100";
        when 9422 => y_in <= "10100100"; x_in <= "01001110"; z_correct<="1110001111111000";
        when 9423 => y_in <= "10100100"; x_in <= "01001111"; z_correct<="1110001110011100";
        when 9424 => y_in <= "10100100"; x_in <= "01010000"; z_correct<="1110001101000000";
        when 9425 => y_in <= "10100100"; x_in <= "01010001"; z_correct<="1110001011100100";
        when 9426 => y_in <= "10100100"; x_in <= "01010010"; z_correct<="1110001010001000";
        when 9427 => y_in <= "10100100"; x_in <= "01010011"; z_correct<="1110001000101100";
        when 9428 => y_in <= "10100100"; x_in <= "01010100"; z_correct<="1110000111010000";
        when 9429 => y_in <= "10100100"; x_in <= "01010101"; z_correct<="1110000101110100";
        when 9430 => y_in <= "10100100"; x_in <= "01010110"; z_correct<="1110000100011000";
        when 9431 => y_in <= "10100100"; x_in <= "01010111"; z_correct<="1110000010111100";
        when 9432 => y_in <= "10100100"; x_in <= "01011000"; z_correct<="1110000001100000";
        when 9433 => y_in <= "10100100"; x_in <= "01011001"; z_correct<="1110000000000100";
        when 9434 => y_in <= "10100100"; x_in <= "01011010"; z_correct<="1101111110101000";
        when 9435 => y_in <= "10100100"; x_in <= "01011011"; z_correct<="1101111101001100";
        when 9436 => y_in <= "10100100"; x_in <= "01011100"; z_correct<="1101111011110000";
        when 9437 => y_in <= "10100100"; x_in <= "01011101"; z_correct<="1101111010010100";
        when 9438 => y_in <= "10100100"; x_in <= "01011110"; z_correct<="1101111000111000";
        when 9439 => y_in <= "10100100"; x_in <= "01011111"; z_correct<="1101110111011100";
        when 9440 => y_in <= "10100100"; x_in <= "01100000"; z_correct<="1101110110000000";
        when 9441 => y_in <= "10100100"; x_in <= "01100001"; z_correct<="1101110100100100";
        when 9442 => y_in <= "10100100"; x_in <= "01100010"; z_correct<="1101110011001000";
        when 9443 => y_in <= "10100100"; x_in <= "01100011"; z_correct<="1101110001101100";
        when 9444 => y_in <= "10100100"; x_in <= "01100100"; z_correct<="1101110000010000";
        when 9445 => y_in <= "10100100"; x_in <= "01100101"; z_correct<="1101101110110100";
        when 9446 => y_in <= "10100100"; x_in <= "01100110"; z_correct<="1101101101011000";
        when 9447 => y_in <= "10100100"; x_in <= "01100111"; z_correct<="1101101011111100";
        when 9448 => y_in <= "10100100"; x_in <= "01101000"; z_correct<="1101101010100000";
        when 9449 => y_in <= "10100100"; x_in <= "01101001"; z_correct<="1101101001000100";
        when 9450 => y_in <= "10100100"; x_in <= "01101010"; z_correct<="1101100111101000";
        when 9451 => y_in <= "10100100"; x_in <= "01101011"; z_correct<="1101100110001100";
        when 9452 => y_in <= "10100100"; x_in <= "01101100"; z_correct<="1101100100110000";
        when 9453 => y_in <= "10100100"; x_in <= "01101101"; z_correct<="1101100011010100";
        when 9454 => y_in <= "10100100"; x_in <= "01101110"; z_correct<="1101100001111000";
        when 9455 => y_in <= "10100100"; x_in <= "01101111"; z_correct<="1101100000011100";
        when 9456 => y_in <= "10100100"; x_in <= "01110000"; z_correct<="1101011111000000";
        when 9457 => y_in <= "10100100"; x_in <= "01110001"; z_correct<="1101011101100100";
        when 9458 => y_in <= "10100100"; x_in <= "01110010"; z_correct<="1101011100001000";
        when 9459 => y_in <= "10100100"; x_in <= "01110011"; z_correct<="1101011010101100";
        when 9460 => y_in <= "10100100"; x_in <= "01110100"; z_correct<="1101011001010000";
        when 9461 => y_in <= "10100100"; x_in <= "01110101"; z_correct<="1101010111110100";
        when 9462 => y_in <= "10100100"; x_in <= "01110110"; z_correct<="1101010110011000";
        when 9463 => y_in <= "10100100"; x_in <= "01110111"; z_correct<="1101010100111100";
        when 9464 => y_in <= "10100100"; x_in <= "01111000"; z_correct<="1101010011100000";
        when 9465 => y_in <= "10100100"; x_in <= "01111001"; z_correct<="1101010010000100";
        when 9466 => y_in <= "10100100"; x_in <= "01111010"; z_correct<="1101010000101000";
        when 9467 => y_in <= "10100100"; x_in <= "01111011"; z_correct<="1101001111001100";
        when 9468 => y_in <= "10100100"; x_in <= "01111100"; z_correct<="1101001101110000";
        when 9469 => y_in <= "10100100"; x_in <= "01111101"; z_correct<="1101001100010100";
        when 9470 => y_in <= "10100100"; x_in <= "01111110"; z_correct<="1101001010111000";
        when 9471 => y_in <= "10100100"; x_in <= "01111111"; z_correct<="1101001001011100";
        when 9472 => y_in <= "10100101"; x_in <= "10000000"; z_correct<="0010110110000000";
        when 9473 => y_in <= "10100101"; x_in <= "10000001"; z_correct<="0010110100100101";
        when 9474 => y_in <= "10100101"; x_in <= "10000010"; z_correct<="0010110011001010";
        when 9475 => y_in <= "10100101"; x_in <= "10000011"; z_correct<="0010110001101111";
        when 9476 => y_in <= "10100101"; x_in <= "10000100"; z_correct<="0010110000010100";
        when 9477 => y_in <= "10100101"; x_in <= "10000101"; z_correct<="0010101110111001";
        when 9478 => y_in <= "10100101"; x_in <= "10000110"; z_correct<="0010101101011110";
        when 9479 => y_in <= "10100101"; x_in <= "10000111"; z_correct<="0010101100000011";
        when 9480 => y_in <= "10100101"; x_in <= "10001000"; z_correct<="0010101010101000";
        when 9481 => y_in <= "10100101"; x_in <= "10001001"; z_correct<="0010101001001101";
        when 9482 => y_in <= "10100101"; x_in <= "10001010"; z_correct<="0010100111110010";
        when 9483 => y_in <= "10100101"; x_in <= "10001011"; z_correct<="0010100110010111";
        when 9484 => y_in <= "10100101"; x_in <= "10001100"; z_correct<="0010100100111100";
        when 9485 => y_in <= "10100101"; x_in <= "10001101"; z_correct<="0010100011100001";
        when 9486 => y_in <= "10100101"; x_in <= "10001110"; z_correct<="0010100010000110";
        when 9487 => y_in <= "10100101"; x_in <= "10001111"; z_correct<="0010100000101011";
        when 9488 => y_in <= "10100101"; x_in <= "10010000"; z_correct<="0010011111010000";
        when 9489 => y_in <= "10100101"; x_in <= "10010001"; z_correct<="0010011101110101";
        when 9490 => y_in <= "10100101"; x_in <= "10010010"; z_correct<="0010011100011010";
        when 9491 => y_in <= "10100101"; x_in <= "10010011"; z_correct<="0010011010111111";
        when 9492 => y_in <= "10100101"; x_in <= "10010100"; z_correct<="0010011001100100";
        when 9493 => y_in <= "10100101"; x_in <= "10010101"; z_correct<="0010011000001001";
        when 9494 => y_in <= "10100101"; x_in <= "10010110"; z_correct<="0010010110101110";
        when 9495 => y_in <= "10100101"; x_in <= "10010111"; z_correct<="0010010101010011";
        when 9496 => y_in <= "10100101"; x_in <= "10011000"; z_correct<="0010010011111000";
        when 9497 => y_in <= "10100101"; x_in <= "10011001"; z_correct<="0010010010011101";
        when 9498 => y_in <= "10100101"; x_in <= "10011010"; z_correct<="0010010001000010";
        when 9499 => y_in <= "10100101"; x_in <= "10011011"; z_correct<="0010001111100111";
        when 9500 => y_in <= "10100101"; x_in <= "10011100"; z_correct<="0010001110001100";
        when 9501 => y_in <= "10100101"; x_in <= "10011101"; z_correct<="0010001100110001";
        when 9502 => y_in <= "10100101"; x_in <= "10011110"; z_correct<="0010001011010110";
        when 9503 => y_in <= "10100101"; x_in <= "10011111"; z_correct<="0010001001111011";
        when 9504 => y_in <= "10100101"; x_in <= "10100000"; z_correct<="0010001000100000";
        when 9505 => y_in <= "10100101"; x_in <= "10100001"; z_correct<="0010000111000101";
        when 9506 => y_in <= "10100101"; x_in <= "10100010"; z_correct<="0010000101101010";
        when 9507 => y_in <= "10100101"; x_in <= "10100011"; z_correct<="0010000100001111";
        when 9508 => y_in <= "10100101"; x_in <= "10100100"; z_correct<="0010000010110100";
        when 9509 => y_in <= "10100101"; x_in <= "10100101"; z_correct<="0010000001011001";
        when 9510 => y_in <= "10100101"; x_in <= "10100110"; z_correct<="0001111111111110";
        when 9511 => y_in <= "10100101"; x_in <= "10100111"; z_correct<="0001111110100011";
        when 9512 => y_in <= "10100101"; x_in <= "10101000"; z_correct<="0001111101001000";
        when 9513 => y_in <= "10100101"; x_in <= "10101001"; z_correct<="0001111011101101";
        when 9514 => y_in <= "10100101"; x_in <= "10101010"; z_correct<="0001111010010010";
        when 9515 => y_in <= "10100101"; x_in <= "10101011"; z_correct<="0001111000110111";
        when 9516 => y_in <= "10100101"; x_in <= "10101100"; z_correct<="0001110111011100";
        when 9517 => y_in <= "10100101"; x_in <= "10101101"; z_correct<="0001110110000001";
        when 9518 => y_in <= "10100101"; x_in <= "10101110"; z_correct<="0001110100100110";
        when 9519 => y_in <= "10100101"; x_in <= "10101111"; z_correct<="0001110011001011";
        when 9520 => y_in <= "10100101"; x_in <= "10110000"; z_correct<="0001110001110000";
        when 9521 => y_in <= "10100101"; x_in <= "10110001"; z_correct<="0001110000010101";
        when 9522 => y_in <= "10100101"; x_in <= "10110010"; z_correct<="0001101110111010";
        when 9523 => y_in <= "10100101"; x_in <= "10110011"; z_correct<="0001101101011111";
        when 9524 => y_in <= "10100101"; x_in <= "10110100"; z_correct<="0001101100000100";
        when 9525 => y_in <= "10100101"; x_in <= "10110101"; z_correct<="0001101010101001";
        when 9526 => y_in <= "10100101"; x_in <= "10110110"; z_correct<="0001101001001110";
        when 9527 => y_in <= "10100101"; x_in <= "10110111"; z_correct<="0001100111110011";
        when 9528 => y_in <= "10100101"; x_in <= "10111000"; z_correct<="0001100110011000";
        when 9529 => y_in <= "10100101"; x_in <= "10111001"; z_correct<="0001100100111101";
        when 9530 => y_in <= "10100101"; x_in <= "10111010"; z_correct<="0001100011100010";
        when 9531 => y_in <= "10100101"; x_in <= "10111011"; z_correct<="0001100010000111";
        when 9532 => y_in <= "10100101"; x_in <= "10111100"; z_correct<="0001100000101100";
        when 9533 => y_in <= "10100101"; x_in <= "10111101"; z_correct<="0001011111010001";
        when 9534 => y_in <= "10100101"; x_in <= "10111110"; z_correct<="0001011101110110";
        when 9535 => y_in <= "10100101"; x_in <= "10111111"; z_correct<="0001011100011011";
        when 9536 => y_in <= "10100101"; x_in <= "11000000"; z_correct<="0001011011000000";
        when 9537 => y_in <= "10100101"; x_in <= "11000001"; z_correct<="0001011001100101";
        when 9538 => y_in <= "10100101"; x_in <= "11000010"; z_correct<="0001011000001010";
        when 9539 => y_in <= "10100101"; x_in <= "11000011"; z_correct<="0001010110101111";
        when 9540 => y_in <= "10100101"; x_in <= "11000100"; z_correct<="0001010101010100";
        when 9541 => y_in <= "10100101"; x_in <= "11000101"; z_correct<="0001010011111001";
        when 9542 => y_in <= "10100101"; x_in <= "11000110"; z_correct<="0001010010011110";
        when 9543 => y_in <= "10100101"; x_in <= "11000111"; z_correct<="0001010001000011";
        when 9544 => y_in <= "10100101"; x_in <= "11001000"; z_correct<="0001001111101000";
        when 9545 => y_in <= "10100101"; x_in <= "11001001"; z_correct<="0001001110001101";
        when 9546 => y_in <= "10100101"; x_in <= "11001010"; z_correct<="0001001100110010";
        when 9547 => y_in <= "10100101"; x_in <= "11001011"; z_correct<="0001001011010111";
        when 9548 => y_in <= "10100101"; x_in <= "11001100"; z_correct<="0001001001111100";
        when 9549 => y_in <= "10100101"; x_in <= "11001101"; z_correct<="0001001000100001";
        when 9550 => y_in <= "10100101"; x_in <= "11001110"; z_correct<="0001000111000110";
        when 9551 => y_in <= "10100101"; x_in <= "11001111"; z_correct<="0001000101101011";
        when 9552 => y_in <= "10100101"; x_in <= "11010000"; z_correct<="0001000100010000";
        when 9553 => y_in <= "10100101"; x_in <= "11010001"; z_correct<="0001000010110101";
        when 9554 => y_in <= "10100101"; x_in <= "11010010"; z_correct<="0001000001011010";
        when 9555 => y_in <= "10100101"; x_in <= "11010011"; z_correct<="0000111111111111";
        when 9556 => y_in <= "10100101"; x_in <= "11010100"; z_correct<="0000111110100100";
        when 9557 => y_in <= "10100101"; x_in <= "11010101"; z_correct<="0000111101001001";
        when 9558 => y_in <= "10100101"; x_in <= "11010110"; z_correct<="0000111011101110";
        when 9559 => y_in <= "10100101"; x_in <= "11010111"; z_correct<="0000111010010011";
        when 9560 => y_in <= "10100101"; x_in <= "11011000"; z_correct<="0000111000111000";
        when 9561 => y_in <= "10100101"; x_in <= "11011001"; z_correct<="0000110111011101";
        when 9562 => y_in <= "10100101"; x_in <= "11011010"; z_correct<="0000110110000010";
        when 9563 => y_in <= "10100101"; x_in <= "11011011"; z_correct<="0000110100100111";
        when 9564 => y_in <= "10100101"; x_in <= "11011100"; z_correct<="0000110011001100";
        when 9565 => y_in <= "10100101"; x_in <= "11011101"; z_correct<="0000110001110001";
        when 9566 => y_in <= "10100101"; x_in <= "11011110"; z_correct<="0000110000010110";
        when 9567 => y_in <= "10100101"; x_in <= "11011111"; z_correct<="0000101110111011";
        when 9568 => y_in <= "10100101"; x_in <= "11100000"; z_correct<="0000101101100000";
        when 9569 => y_in <= "10100101"; x_in <= "11100001"; z_correct<="0000101100000101";
        when 9570 => y_in <= "10100101"; x_in <= "11100010"; z_correct<="0000101010101010";
        when 9571 => y_in <= "10100101"; x_in <= "11100011"; z_correct<="0000101001001111";
        when 9572 => y_in <= "10100101"; x_in <= "11100100"; z_correct<="0000100111110100";
        when 9573 => y_in <= "10100101"; x_in <= "11100101"; z_correct<="0000100110011001";
        when 9574 => y_in <= "10100101"; x_in <= "11100110"; z_correct<="0000100100111110";
        when 9575 => y_in <= "10100101"; x_in <= "11100111"; z_correct<="0000100011100011";
        when 9576 => y_in <= "10100101"; x_in <= "11101000"; z_correct<="0000100010001000";
        when 9577 => y_in <= "10100101"; x_in <= "11101001"; z_correct<="0000100000101101";
        when 9578 => y_in <= "10100101"; x_in <= "11101010"; z_correct<="0000011111010010";
        when 9579 => y_in <= "10100101"; x_in <= "11101011"; z_correct<="0000011101110111";
        when 9580 => y_in <= "10100101"; x_in <= "11101100"; z_correct<="0000011100011100";
        when 9581 => y_in <= "10100101"; x_in <= "11101101"; z_correct<="0000011011000001";
        when 9582 => y_in <= "10100101"; x_in <= "11101110"; z_correct<="0000011001100110";
        when 9583 => y_in <= "10100101"; x_in <= "11101111"; z_correct<="0000011000001011";
        when 9584 => y_in <= "10100101"; x_in <= "11110000"; z_correct<="0000010110110000";
        when 9585 => y_in <= "10100101"; x_in <= "11110001"; z_correct<="0000010101010101";
        when 9586 => y_in <= "10100101"; x_in <= "11110010"; z_correct<="0000010011111010";
        when 9587 => y_in <= "10100101"; x_in <= "11110011"; z_correct<="0000010010011111";
        when 9588 => y_in <= "10100101"; x_in <= "11110100"; z_correct<="0000010001000100";
        when 9589 => y_in <= "10100101"; x_in <= "11110101"; z_correct<="0000001111101001";
        when 9590 => y_in <= "10100101"; x_in <= "11110110"; z_correct<="0000001110001110";
        when 9591 => y_in <= "10100101"; x_in <= "11110111"; z_correct<="0000001100110011";
        when 9592 => y_in <= "10100101"; x_in <= "11111000"; z_correct<="0000001011011000";
        when 9593 => y_in <= "10100101"; x_in <= "11111001"; z_correct<="0000001001111101";
        when 9594 => y_in <= "10100101"; x_in <= "11111010"; z_correct<="0000001000100010";
        when 9595 => y_in <= "10100101"; x_in <= "11111011"; z_correct<="0000000111000111";
        when 9596 => y_in <= "10100101"; x_in <= "11111100"; z_correct<="0000000101101100";
        when 9597 => y_in <= "10100101"; x_in <= "11111101"; z_correct<="0000000100010001";
        when 9598 => y_in <= "10100101"; x_in <= "11111110"; z_correct<="0000000010110110";
        when 9599 => y_in <= "10100101"; x_in <= "11111111"; z_correct<="0000000001011011";
        when 9600 => y_in <= "10100101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 9601 => y_in <= "10100101"; x_in <= "00000001"; z_correct<="1111111110100101";
        when 9602 => y_in <= "10100101"; x_in <= "00000010"; z_correct<="1111111101001010";
        when 9603 => y_in <= "10100101"; x_in <= "00000011"; z_correct<="1111111011101111";
        when 9604 => y_in <= "10100101"; x_in <= "00000100"; z_correct<="1111111010010100";
        when 9605 => y_in <= "10100101"; x_in <= "00000101"; z_correct<="1111111000111001";
        when 9606 => y_in <= "10100101"; x_in <= "00000110"; z_correct<="1111110111011110";
        when 9607 => y_in <= "10100101"; x_in <= "00000111"; z_correct<="1111110110000011";
        when 9608 => y_in <= "10100101"; x_in <= "00001000"; z_correct<="1111110100101000";
        when 9609 => y_in <= "10100101"; x_in <= "00001001"; z_correct<="1111110011001101";
        when 9610 => y_in <= "10100101"; x_in <= "00001010"; z_correct<="1111110001110010";
        when 9611 => y_in <= "10100101"; x_in <= "00001011"; z_correct<="1111110000010111";
        when 9612 => y_in <= "10100101"; x_in <= "00001100"; z_correct<="1111101110111100";
        when 9613 => y_in <= "10100101"; x_in <= "00001101"; z_correct<="1111101101100001";
        when 9614 => y_in <= "10100101"; x_in <= "00001110"; z_correct<="1111101100000110";
        when 9615 => y_in <= "10100101"; x_in <= "00001111"; z_correct<="1111101010101011";
        when 9616 => y_in <= "10100101"; x_in <= "00010000"; z_correct<="1111101001010000";
        when 9617 => y_in <= "10100101"; x_in <= "00010001"; z_correct<="1111100111110101";
        when 9618 => y_in <= "10100101"; x_in <= "00010010"; z_correct<="1111100110011010";
        when 9619 => y_in <= "10100101"; x_in <= "00010011"; z_correct<="1111100100111111";
        when 9620 => y_in <= "10100101"; x_in <= "00010100"; z_correct<="1111100011100100";
        when 9621 => y_in <= "10100101"; x_in <= "00010101"; z_correct<="1111100010001001";
        when 9622 => y_in <= "10100101"; x_in <= "00010110"; z_correct<="1111100000101110";
        when 9623 => y_in <= "10100101"; x_in <= "00010111"; z_correct<="1111011111010011";
        when 9624 => y_in <= "10100101"; x_in <= "00011000"; z_correct<="1111011101111000";
        when 9625 => y_in <= "10100101"; x_in <= "00011001"; z_correct<="1111011100011101";
        when 9626 => y_in <= "10100101"; x_in <= "00011010"; z_correct<="1111011011000010";
        when 9627 => y_in <= "10100101"; x_in <= "00011011"; z_correct<="1111011001100111";
        when 9628 => y_in <= "10100101"; x_in <= "00011100"; z_correct<="1111011000001100";
        when 9629 => y_in <= "10100101"; x_in <= "00011101"; z_correct<="1111010110110001";
        when 9630 => y_in <= "10100101"; x_in <= "00011110"; z_correct<="1111010101010110";
        when 9631 => y_in <= "10100101"; x_in <= "00011111"; z_correct<="1111010011111011";
        when 9632 => y_in <= "10100101"; x_in <= "00100000"; z_correct<="1111010010100000";
        when 9633 => y_in <= "10100101"; x_in <= "00100001"; z_correct<="1111010001000101";
        when 9634 => y_in <= "10100101"; x_in <= "00100010"; z_correct<="1111001111101010";
        when 9635 => y_in <= "10100101"; x_in <= "00100011"; z_correct<="1111001110001111";
        when 9636 => y_in <= "10100101"; x_in <= "00100100"; z_correct<="1111001100110100";
        when 9637 => y_in <= "10100101"; x_in <= "00100101"; z_correct<="1111001011011001";
        when 9638 => y_in <= "10100101"; x_in <= "00100110"; z_correct<="1111001001111110";
        when 9639 => y_in <= "10100101"; x_in <= "00100111"; z_correct<="1111001000100011";
        when 9640 => y_in <= "10100101"; x_in <= "00101000"; z_correct<="1111000111001000";
        when 9641 => y_in <= "10100101"; x_in <= "00101001"; z_correct<="1111000101101101";
        when 9642 => y_in <= "10100101"; x_in <= "00101010"; z_correct<="1111000100010010";
        when 9643 => y_in <= "10100101"; x_in <= "00101011"; z_correct<="1111000010110111";
        when 9644 => y_in <= "10100101"; x_in <= "00101100"; z_correct<="1111000001011100";
        when 9645 => y_in <= "10100101"; x_in <= "00101101"; z_correct<="1111000000000001";
        when 9646 => y_in <= "10100101"; x_in <= "00101110"; z_correct<="1110111110100110";
        when 9647 => y_in <= "10100101"; x_in <= "00101111"; z_correct<="1110111101001011";
        when 9648 => y_in <= "10100101"; x_in <= "00110000"; z_correct<="1110111011110000";
        when 9649 => y_in <= "10100101"; x_in <= "00110001"; z_correct<="1110111010010101";
        when 9650 => y_in <= "10100101"; x_in <= "00110010"; z_correct<="1110111000111010";
        when 9651 => y_in <= "10100101"; x_in <= "00110011"; z_correct<="1110110111011111";
        when 9652 => y_in <= "10100101"; x_in <= "00110100"; z_correct<="1110110110000100";
        when 9653 => y_in <= "10100101"; x_in <= "00110101"; z_correct<="1110110100101001";
        when 9654 => y_in <= "10100101"; x_in <= "00110110"; z_correct<="1110110011001110";
        when 9655 => y_in <= "10100101"; x_in <= "00110111"; z_correct<="1110110001110011";
        when 9656 => y_in <= "10100101"; x_in <= "00111000"; z_correct<="1110110000011000";
        when 9657 => y_in <= "10100101"; x_in <= "00111001"; z_correct<="1110101110111101";
        when 9658 => y_in <= "10100101"; x_in <= "00111010"; z_correct<="1110101101100010";
        when 9659 => y_in <= "10100101"; x_in <= "00111011"; z_correct<="1110101100000111";
        when 9660 => y_in <= "10100101"; x_in <= "00111100"; z_correct<="1110101010101100";
        when 9661 => y_in <= "10100101"; x_in <= "00111101"; z_correct<="1110101001010001";
        when 9662 => y_in <= "10100101"; x_in <= "00111110"; z_correct<="1110100111110110";
        when 9663 => y_in <= "10100101"; x_in <= "00111111"; z_correct<="1110100110011011";
        when 9664 => y_in <= "10100101"; x_in <= "01000000"; z_correct<="1110100101000000";
        when 9665 => y_in <= "10100101"; x_in <= "01000001"; z_correct<="1110100011100101";
        when 9666 => y_in <= "10100101"; x_in <= "01000010"; z_correct<="1110100010001010";
        when 9667 => y_in <= "10100101"; x_in <= "01000011"; z_correct<="1110100000101111";
        when 9668 => y_in <= "10100101"; x_in <= "01000100"; z_correct<="1110011111010100";
        when 9669 => y_in <= "10100101"; x_in <= "01000101"; z_correct<="1110011101111001";
        when 9670 => y_in <= "10100101"; x_in <= "01000110"; z_correct<="1110011100011110";
        when 9671 => y_in <= "10100101"; x_in <= "01000111"; z_correct<="1110011011000011";
        when 9672 => y_in <= "10100101"; x_in <= "01001000"; z_correct<="1110011001101000";
        when 9673 => y_in <= "10100101"; x_in <= "01001001"; z_correct<="1110011000001101";
        when 9674 => y_in <= "10100101"; x_in <= "01001010"; z_correct<="1110010110110010";
        when 9675 => y_in <= "10100101"; x_in <= "01001011"; z_correct<="1110010101010111";
        when 9676 => y_in <= "10100101"; x_in <= "01001100"; z_correct<="1110010011111100";
        when 9677 => y_in <= "10100101"; x_in <= "01001101"; z_correct<="1110010010100001";
        when 9678 => y_in <= "10100101"; x_in <= "01001110"; z_correct<="1110010001000110";
        when 9679 => y_in <= "10100101"; x_in <= "01001111"; z_correct<="1110001111101011";
        when 9680 => y_in <= "10100101"; x_in <= "01010000"; z_correct<="1110001110010000";
        when 9681 => y_in <= "10100101"; x_in <= "01010001"; z_correct<="1110001100110101";
        when 9682 => y_in <= "10100101"; x_in <= "01010010"; z_correct<="1110001011011010";
        when 9683 => y_in <= "10100101"; x_in <= "01010011"; z_correct<="1110001001111111";
        when 9684 => y_in <= "10100101"; x_in <= "01010100"; z_correct<="1110001000100100";
        when 9685 => y_in <= "10100101"; x_in <= "01010101"; z_correct<="1110000111001001";
        when 9686 => y_in <= "10100101"; x_in <= "01010110"; z_correct<="1110000101101110";
        when 9687 => y_in <= "10100101"; x_in <= "01010111"; z_correct<="1110000100010011";
        when 9688 => y_in <= "10100101"; x_in <= "01011000"; z_correct<="1110000010111000";
        when 9689 => y_in <= "10100101"; x_in <= "01011001"; z_correct<="1110000001011101";
        when 9690 => y_in <= "10100101"; x_in <= "01011010"; z_correct<="1110000000000010";
        when 9691 => y_in <= "10100101"; x_in <= "01011011"; z_correct<="1101111110100111";
        when 9692 => y_in <= "10100101"; x_in <= "01011100"; z_correct<="1101111101001100";
        when 9693 => y_in <= "10100101"; x_in <= "01011101"; z_correct<="1101111011110001";
        when 9694 => y_in <= "10100101"; x_in <= "01011110"; z_correct<="1101111010010110";
        when 9695 => y_in <= "10100101"; x_in <= "01011111"; z_correct<="1101111000111011";
        when 9696 => y_in <= "10100101"; x_in <= "01100000"; z_correct<="1101110111100000";
        when 9697 => y_in <= "10100101"; x_in <= "01100001"; z_correct<="1101110110000101";
        when 9698 => y_in <= "10100101"; x_in <= "01100010"; z_correct<="1101110100101010";
        when 9699 => y_in <= "10100101"; x_in <= "01100011"; z_correct<="1101110011001111";
        when 9700 => y_in <= "10100101"; x_in <= "01100100"; z_correct<="1101110001110100";
        when 9701 => y_in <= "10100101"; x_in <= "01100101"; z_correct<="1101110000011001";
        when 9702 => y_in <= "10100101"; x_in <= "01100110"; z_correct<="1101101110111110";
        when 9703 => y_in <= "10100101"; x_in <= "01100111"; z_correct<="1101101101100011";
        when 9704 => y_in <= "10100101"; x_in <= "01101000"; z_correct<="1101101100001000";
        when 9705 => y_in <= "10100101"; x_in <= "01101001"; z_correct<="1101101010101101";
        when 9706 => y_in <= "10100101"; x_in <= "01101010"; z_correct<="1101101001010010";
        when 9707 => y_in <= "10100101"; x_in <= "01101011"; z_correct<="1101100111110111";
        when 9708 => y_in <= "10100101"; x_in <= "01101100"; z_correct<="1101100110011100";
        when 9709 => y_in <= "10100101"; x_in <= "01101101"; z_correct<="1101100101000001";
        when 9710 => y_in <= "10100101"; x_in <= "01101110"; z_correct<="1101100011100110";
        when 9711 => y_in <= "10100101"; x_in <= "01101111"; z_correct<="1101100010001011";
        when 9712 => y_in <= "10100101"; x_in <= "01110000"; z_correct<="1101100000110000";
        when 9713 => y_in <= "10100101"; x_in <= "01110001"; z_correct<="1101011111010101";
        when 9714 => y_in <= "10100101"; x_in <= "01110010"; z_correct<="1101011101111010";
        when 9715 => y_in <= "10100101"; x_in <= "01110011"; z_correct<="1101011100011111";
        when 9716 => y_in <= "10100101"; x_in <= "01110100"; z_correct<="1101011011000100";
        when 9717 => y_in <= "10100101"; x_in <= "01110101"; z_correct<="1101011001101001";
        when 9718 => y_in <= "10100101"; x_in <= "01110110"; z_correct<="1101011000001110";
        when 9719 => y_in <= "10100101"; x_in <= "01110111"; z_correct<="1101010110110011";
        when 9720 => y_in <= "10100101"; x_in <= "01111000"; z_correct<="1101010101011000";
        when 9721 => y_in <= "10100101"; x_in <= "01111001"; z_correct<="1101010011111101";
        when 9722 => y_in <= "10100101"; x_in <= "01111010"; z_correct<="1101010010100010";
        when 9723 => y_in <= "10100101"; x_in <= "01111011"; z_correct<="1101010001000111";
        when 9724 => y_in <= "10100101"; x_in <= "01111100"; z_correct<="1101001111101100";
        when 9725 => y_in <= "10100101"; x_in <= "01111101"; z_correct<="1101001110010001";
        when 9726 => y_in <= "10100101"; x_in <= "01111110"; z_correct<="1101001100110110";
        when 9727 => y_in <= "10100101"; x_in <= "01111111"; z_correct<="1101001011011011";
        when 9728 => y_in <= "10100110"; x_in <= "10000000"; z_correct<="0010110100000000";
        when 9729 => y_in <= "10100110"; x_in <= "10000001"; z_correct<="0010110010100110";
        when 9730 => y_in <= "10100110"; x_in <= "10000010"; z_correct<="0010110001001100";
        when 9731 => y_in <= "10100110"; x_in <= "10000011"; z_correct<="0010101111110010";
        when 9732 => y_in <= "10100110"; x_in <= "10000100"; z_correct<="0010101110011000";
        when 9733 => y_in <= "10100110"; x_in <= "10000101"; z_correct<="0010101100111110";
        when 9734 => y_in <= "10100110"; x_in <= "10000110"; z_correct<="0010101011100100";
        when 9735 => y_in <= "10100110"; x_in <= "10000111"; z_correct<="0010101010001010";
        when 9736 => y_in <= "10100110"; x_in <= "10001000"; z_correct<="0010101000110000";
        when 9737 => y_in <= "10100110"; x_in <= "10001001"; z_correct<="0010100111010110";
        when 9738 => y_in <= "10100110"; x_in <= "10001010"; z_correct<="0010100101111100";
        when 9739 => y_in <= "10100110"; x_in <= "10001011"; z_correct<="0010100100100010";
        when 9740 => y_in <= "10100110"; x_in <= "10001100"; z_correct<="0010100011001000";
        when 9741 => y_in <= "10100110"; x_in <= "10001101"; z_correct<="0010100001101110";
        when 9742 => y_in <= "10100110"; x_in <= "10001110"; z_correct<="0010100000010100";
        when 9743 => y_in <= "10100110"; x_in <= "10001111"; z_correct<="0010011110111010";
        when 9744 => y_in <= "10100110"; x_in <= "10010000"; z_correct<="0010011101100000";
        when 9745 => y_in <= "10100110"; x_in <= "10010001"; z_correct<="0010011100000110";
        when 9746 => y_in <= "10100110"; x_in <= "10010010"; z_correct<="0010011010101100";
        when 9747 => y_in <= "10100110"; x_in <= "10010011"; z_correct<="0010011001010010";
        when 9748 => y_in <= "10100110"; x_in <= "10010100"; z_correct<="0010010111111000";
        when 9749 => y_in <= "10100110"; x_in <= "10010101"; z_correct<="0010010110011110";
        when 9750 => y_in <= "10100110"; x_in <= "10010110"; z_correct<="0010010101000100";
        when 9751 => y_in <= "10100110"; x_in <= "10010111"; z_correct<="0010010011101010";
        when 9752 => y_in <= "10100110"; x_in <= "10011000"; z_correct<="0010010010010000";
        when 9753 => y_in <= "10100110"; x_in <= "10011001"; z_correct<="0010010000110110";
        when 9754 => y_in <= "10100110"; x_in <= "10011010"; z_correct<="0010001111011100";
        when 9755 => y_in <= "10100110"; x_in <= "10011011"; z_correct<="0010001110000010";
        when 9756 => y_in <= "10100110"; x_in <= "10011100"; z_correct<="0010001100101000";
        when 9757 => y_in <= "10100110"; x_in <= "10011101"; z_correct<="0010001011001110";
        when 9758 => y_in <= "10100110"; x_in <= "10011110"; z_correct<="0010001001110100";
        when 9759 => y_in <= "10100110"; x_in <= "10011111"; z_correct<="0010001000011010";
        when 9760 => y_in <= "10100110"; x_in <= "10100000"; z_correct<="0010000111000000";
        when 9761 => y_in <= "10100110"; x_in <= "10100001"; z_correct<="0010000101100110";
        when 9762 => y_in <= "10100110"; x_in <= "10100010"; z_correct<="0010000100001100";
        when 9763 => y_in <= "10100110"; x_in <= "10100011"; z_correct<="0010000010110010";
        when 9764 => y_in <= "10100110"; x_in <= "10100100"; z_correct<="0010000001011000";
        when 9765 => y_in <= "10100110"; x_in <= "10100101"; z_correct<="0001111111111110";
        when 9766 => y_in <= "10100110"; x_in <= "10100110"; z_correct<="0001111110100100";
        when 9767 => y_in <= "10100110"; x_in <= "10100111"; z_correct<="0001111101001010";
        when 9768 => y_in <= "10100110"; x_in <= "10101000"; z_correct<="0001111011110000";
        when 9769 => y_in <= "10100110"; x_in <= "10101001"; z_correct<="0001111010010110";
        when 9770 => y_in <= "10100110"; x_in <= "10101010"; z_correct<="0001111000111100";
        when 9771 => y_in <= "10100110"; x_in <= "10101011"; z_correct<="0001110111100010";
        when 9772 => y_in <= "10100110"; x_in <= "10101100"; z_correct<="0001110110001000";
        when 9773 => y_in <= "10100110"; x_in <= "10101101"; z_correct<="0001110100101110";
        when 9774 => y_in <= "10100110"; x_in <= "10101110"; z_correct<="0001110011010100";
        when 9775 => y_in <= "10100110"; x_in <= "10101111"; z_correct<="0001110001111010";
        when 9776 => y_in <= "10100110"; x_in <= "10110000"; z_correct<="0001110000100000";
        when 9777 => y_in <= "10100110"; x_in <= "10110001"; z_correct<="0001101111000110";
        when 9778 => y_in <= "10100110"; x_in <= "10110010"; z_correct<="0001101101101100";
        when 9779 => y_in <= "10100110"; x_in <= "10110011"; z_correct<="0001101100010010";
        when 9780 => y_in <= "10100110"; x_in <= "10110100"; z_correct<="0001101010111000";
        when 9781 => y_in <= "10100110"; x_in <= "10110101"; z_correct<="0001101001011110";
        when 9782 => y_in <= "10100110"; x_in <= "10110110"; z_correct<="0001101000000100";
        when 9783 => y_in <= "10100110"; x_in <= "10110111"; z_correct<="0001100110101010";
        when 9784 => y_in <= "10100110"; x_in <= "10111000"; z_correct<="0001100101010000";
        when 9785 => y_in <= "10100110"; x_in <= "10111001"; z_correct<="0001100011110110";
        when 9786 => y_in <= "10100110"; x_in <= "10111010"; z_correct<="0001100010011100";
        when 9787 => y_in <= "10100110"; x_in <= "10111011"; z_correct<="0001100001000010";
        when 9788 => y_in <= "10100110"; x_in <= "10111100"; z_correct<="0001011111101000";
        when 9789 => y_in <= "10100110"; x_in <= "10111101"; z_correct<="0001011110001110";
        when 9790 => y_in <= "10100110"; x_in <= "10111110"; z_correct<="0001011100110100";
        when 9791 => y_in <= "10100110"; x_in <= "10111111"; z_correct<="0001011011011010";
        when 9792 => y_in <= "10100110"; x_in <= "11000000"; z_correct<="0001011010000000";
        when 9793 => y_in <= "10100110"; x_in <= "11000001"; z_correct<="0001011000100110";
        when 9794 => y_in <= "10100110"; x_in <= "11000010"; z_correct<="0001010111001100";
        when 9795 => y_in <= "10100110"; x_in <= "11000011"; z_correct<="0001010101110010";
        when 9796 => y_in <= "10100110"; x_in <= "11000100"; z_correct<="0001010100011000";
        when 9797 => y_in <= "10100110"; x_in <= "11000101"; z_correct<="0001010010111110";
        when 9798 => y_in <= "10100110"; x_in <= "11000110"; z_correct<="0001010001100100";
        when 9799 => y_in <= "10100110"; x_in <= "11000111"; z_correct<="0001010000001010";
        when 9800 => y_in <= "10100110"; x_in <= "11001000"; z_correct<="0001001110110000";
        when 9801 => y_in <= "10100110"; x_in <= "11001001"; z_correct<="0001001101010110";
        when 9802 => y_in <= "10100110"; x_in <= "11001010"; z_correct<="0001001011111100";
        when 9803 => y_in <= "10100110"; x_in <= "11001011"; z_correct<="0001001010100010";
        when 9804 => y_in <= "10100110"; x_in <= "11001100"; z_correct<="0001001001001000";
        when 9805 => y_in <= "10100110"; x_in <= "11001101"; z_correct<="0001000111101110";
        when 9806 => y_in <= "10100110"; x_in <= "11001110"; z_correct<="0001000110010100";
        when 9807 => y_in <= "10100110"; x_in <= "11001111"; z_correct<="0001000100111010";
        when 9808 => y_in <= "10100110"; x_in <= "11010000"; z_correct<="0001000011100000";
        when 9809 => y_in <= "10100110"; x_in <= "11010001"; z_correct<="0001000010000110";
        when 9810 => y_in <= "10100110"; x_in <= "11010010"; z_correct<="0001000000101100";
        when 9811 => y_in <= "10100110"; x_in <= "11010011"; z_correct<="0000111111010010";
        when 9812 => y_in <= "10100110"; x_in <= "11010100"; z_correct<="0000111101111000";
        when 9813 => y_in <= "10100110"; x_in <= "11010101"; z_correct<="0000111100011110";
        when 9814 => y_in <= "10100110"; x_in <= "11010110"; z_correct<="0000111011000100";
        when 9815 => y_in <= "10100110"; x_in <= "11010111"; z_correct<="0000111001101010";
        when 9816 => y_in <= "10100110"; x_in <= "11011000"; z_correct<="0000111000010000";
        when 9817 => y_in <= "10100110"; x_in <= "11011001"; z_correct<="0000110110110110";
        when 9818 => y_in <= "10100110"; x_in <= "11011010"; z_correct<="0000110101011100";
        when 9819 => y_in <= "10100110"; x_in <= "11011011"; z_correct<="0000110100000010";
        when 9820 => y_in <= "10100110"; x_in <= "11011100"; z_correct<="0000110010101000";
        when 9821 => y_in <= "10100110"; x_in <= "11011101"; z_correct<="0000110001001110";
        when 9822 => y_in <= "10100110"; x_in <= "11011110"; z_correct<="0000101111110100";
        when 9823 => y_in <= "10100110"; x_in <= "11011111"; z_correct<="0000101110011010";
        when 9824 => y_in <= "10100110"; x_in <= "11100000"; z_correct<="0000101101000000";
        when 9825 => y_in <= "10100110"; x_in <= "11100001"; z_correct<="0000101011100110";
        when 9826 => y_in <= "10100110"; x_in <= "11100010"; z_correct<="0000101010001100";
        when 9827 => y_in <= "10100110"; x_in <= "11100011"; z_correct<="0000101000110010";
        when 9828 => y_in <= "10100110"; x_in <= "11100100"; z_correct<="0000100111011000";
        when 9829 => y_in <= "10100110"; x_in <= "11100101"; z_correct<="0000100101111110";
        when 9830 => y_in <= "10100110"; x_in <= "11100110"; z_correct<="0000100100100100";
        when 9831 => y_in <= "10100110"; x_in <= "11100111"; z_correct<="0000100011001010";
        when 9832 => y_in <= "10100110"; x_in <= "11101000"; z_correct<="0000100001110000";
        when 9833 => y_in <= "10100110"; x_in <= "11101001"; z_correct<="0000100000010110";
        when 9834 => y_in <= "10100110"; x_in <= "11101010"; z_correct<="0000011110111100";
        when 9835 => y_in <= "10100110"; x_in <= "11101011"; z_correct<="0000011101100010";
        when 9836 => y_in <= "10100110"; x_in <= "11101100"; z_correct<="0000011100001000";
        when 9837 => y_in <= "10100110"; x_in <= "11101101"; z_correct<="0000011010101110";
        when 9838 => y_in <= "10100110"; x_in <= "11101110"; z_correct<="0000011001010100";
        when 9839 => y_in <= "10100110"; x_in <= "11101111"; z_correct<="0000010111111010";
        when 9840 => y_in <= "10100110"; x_in <= "11110000"; z_correct<="0000010110100000";
        when 9841 => y_in <= "10100110"; x_in <= "11110001"; z_correct<="0000010101000110";
        when 9842 => y_in <= "10100110"; x_in <= "11110010"; z_correct<="0000010011101100";
        when 9843 => y_in <= "10100110"; x_in <= "11110011"; z_correct<="0000010010010010";
        when 9844 => y_in <= "10100110"; x_in <= "11110100"; z_correct<="0000010000111000";
        when 9845 => y_in <= "10100110"; x_in <= "11110101"; z_correct<="0000001111011110";
        when 9846 => y_in <= "10100110"; x_in <= "11110110"; z_correct<="0000001110000100";
        when 9847 => y_in <= "10100110"; x_in <= "11110111"; z_correct<="0000001100101010";
        when 9848 => y_in <= "10100110"; x_in <= "11111000"; z_correct<="0000001011010000";
        when 9849 => y_in <= "10100110"; x_in <= "11111001"; z_correct<="0000001001110110";
        when 9850 => y_in <= "10100110"; x_in <= "11111010"; z_correct<="0000001000011100";
        when 9851 => y_in <= "10100110"; x_in <= "11111011"; z_correct<="0000000111000010";
        when 9852 => y_in <= "10100110"; x_in <= "11111100"; z_correct<="0000000101101000";
        when 9853 => y_in <= "10100110"; x_in <= "11111101"; z_correct<="0000000100001110";
        when 9854 => y_in <= "10100110"; x_in <= "11111110"; z_correct<="0000000010110100";
        when 9855 => y_in <= "10100110"; x_in <= "11111111"; z_correct<="0000000001011010";
        when 9856 => y_in <= "10100110"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 9857 => y_in <= "10100110"; x_in <= "00000001"; z_correct<="1111111110100110";
        when 9858 => y_in <= "10100110"; x_in <= "00000010"; z_correct<="1111111101001100";
        when 9859 => y_in <= "10100110"; x_in <= "00000011"; z_correct<="1111111011110010";
        when 9860 => y_in <= "10100110"; x_in <= "00000100"; z_correct<="1111111010011000";
        when 9861 => y_in <= "10100110"; x_in <= "00000101"; z_correct<="1111111000111110";
        when 9862 => y_in <= "10100110"; x_in <= "00000110"; z_correct<="1111110111100100";
        when 9863 => y_in <= "10100110"; x_in <= "00000111"; z_correct<="1111110110001010";
        when 9864 => y_in <= "10100110"; x_in <= "00001000"; z_correct<="1111110100110000";
        when 9865 => y_in <= "10100110"; x_in <= "00001001"; z_correct<="1111110011010110";
        when 9866 => y_in <= "10100110"; x_in <= "00001010"; z_correct<="1111110001111100";
        when 9867 => y_in <= "10100110"; x_in <= "00001011"; z_correct<="1111110000100010";
        when 9868 => y_in <= "10100110"; x_in <= "00001100"; z_correct<="1111101111001000";
        when 9869 => y_in <= "10100110"; x_in <= "00001101"; z_correct<="1111101101101110";
        when 9870 => y_in <= "10100110"; x_in <= "00001110"; z_correct<="1111101100010100";
        when 9871 => y_in <= "10100110"; x_in <= "00001111"; z_correct<="1111101010111010";
        when 9872 => y_in <= "10100110"; x_in <= "00010000"; z_correct<="1111101001100000";
        when 9873 => y_in <= "10100110"; x_in <= "00010001"; z_correct<="1111101000000110";
        when 9874 => y_in <= "10100110"; x_in <= "00010010"; z_correct<="1111100110101100";
        when 9875 => y_in <= "10100110"; x_in <= "00010011"; z_correct<="1111100101010010";
        when 9876 => y_in <= "10100110"; x_in <= "00010100"; z_correct<="1111100011111000";
        when 9877 => y_in <= "10100110"; x_in <= "00010101"; z_correct<="1111100010011110";
        when 9878 => y_in <= "10100110"; x_in <= "00010110"; z_correct<="1111100001000100";
        when 9879 => y_in <= "10100110"; x_in <= "00010111"; z_correct<="1111011111101010";
        when 9880 => y_in <= "10100110"; x_in <= "00011000"; z_correct<="1111011110010000";
        when 9881 => y_in <= "10100110"; x_in <= "00011001"; z_correct<="1111011100110110";
        when 9882 => y_in <= "10100110"; x_in <= "00011010"; z_correct<="1111011011011100";
        when 9883 => y_in <= "10100110"; x_in <= "00011011"; z_correct<="1111011010000010";
        when 9884 => y_in <= "10100110"; x_in <= "00011100"; z_correct<="1111011000101000";
        when 9885 => y_in <= "10100110"; x_in <= "00011101"; z_correct<="1111010111001110";
        when 9886 => y_in <= "10100110"; x_in <= "00011110"; z_correct<="1111010101110100";
        when 9887 => y_in <= "10100110"; x_in <= "00011111"; z_correct<="1111010100011010";
        when 9888 => y_in <= "10100110"; x_in <= "00100000"; z_correct<="1111010011000000";
        when 9889 => y_in <= "10100110"; x_in <= "00100001"; z_correct<="1111010001100110";
        when 9890 => y_in <= "10100110"; x_in <= "00100010"; z_correct<="1111010000001100";
        when 9891 => y_in <= "10100110"; x_in <= "00100011"; z_correct<="1111001110110010";
        when 9892 => y_in <= "10100110"; x_in <= "00100100"; z_correct<="1111001101011000";
        when 9893 => y_in <= "10100110"; x_in <= "00100101"; z_correct<="1111001011111110";
        when 9894 => y_in <= "10100110"; x_in <= "00100110"; z_correct<="1111001010100100";
        when 9895 => y_in <= "10100110"; x_in <= "00100111"; z_correct<="1111001001001010";
        when 9896 => y_in <= "10100110"; x_in <= "00101000"; z_correct<="1111000111110000";
        when 9897 => y_in <= "10100110"; x_in <= "00101001"; z_correct<="1111000110010110";
        when 9898 => y_in <= "10100110"; x_in <= "00101010"; z_correct<="1111000100111100";
        when 9899 => y_in <= "10100110"; x_in <= "00101011"; z_correct<="1111000011100010";
        when 9900 => y_in <= "10100110"; x_in <= "00101100"; z_correct<="1111000010001000";
        when 9901 => y_in <= "10100110"; x_in <= "00101101"; z_correct<="1111000000101110";
        when 9902 => y_in <= "10100110"; x_in <= "00101110"; z_correct<="1110111111010100";
        when 9903 => y_in <= "10100110"; x_in <= "00101111"; z_correct<="1110111101111010";
        when 9904 => y_in <= "10100110"; x_in <= "00110000"; z_correct<="1110111100100000";
        when 9905 => y_in <= "10100110"; x_in <= "00110001"; z_correct<="1110111011000110";
        when 9906 => y_in <= "10100110"; x_in <= "00110010"; z_correct<="1110111001101100";
        when 9907 => y_in <= "10100110"; x_in <= "00110011"; z_correct<="1110111000010010";
        when 9908 => y_in <= "10100110"; x_in <= "00110100"; z_correct<="1110110110111000";
        when 9909 => y_in <= "10100110"; x_in <= "00110101"; z_correct<="1110110101011110";
        when 9910 => y_in <= "10100110"; x_in <= "00110110"; z_correct<="1110110100000100";
        when 9911 => y_in <= "10100110"; x_in <= "00110111"; z_correct<="1110110010101010";
        when 9912 => y_in <= "10100110"; x_in <= "00111000"; z_correct<="1110110001010000";
        when 9913 => y_in <= "10100110"; x_in <= "00111001"; z_correct<="1110101111110110";
        when 9914 => y_in <= "10100110"; x_in <= "00111010"; z_correct<="1110101110011100";
        when 9915 => y_in <= "10100110"; x_in <= "00111011"; z_correct<="1110101101000010";
        when 9916 => y_in <= "10100110"; x_in <= "00111100"; z_correct<="1110101011101000";
        when 9917 => y_in <= "10100110"; x_in <= "00111101"; z_correct<="1110101010001110";
        when 9918 => y_in <= "10100110"; x_in <= "00111110"; z_correct<="1110101000110100";
        when 9919 => y_in <= "10100110"; x_in <= "00111111"; z_correct<="1110100111011010";
        when 9920 => y_in <= "10100110"; x_in <= "01000000"; z_correct<="1110100110000000";
        when 9921 => y_in <= "10100110"; x_in <= "01000001"; z_correct<="1110100100100110";
        when 9922 => y_in <= "10100110"; x_in <= "01000010"; z_correct<="1110100011001100";
        when 9923 => y_in <= "10100110"; x_in <= "01000011"; z_correct<="1110100001110010";
        when 9924 => y_in <= "10100110"; x_in <= "01000100"; z_correct<="1110100000011000";
        when 9925 => y_in <= "10100110"; x_in <= "01000101"; z_correct<="1110011110111110";
        when 9926 => y_in <= "10100110"; x_in <= "01000110"; z_correct<="1110011101100100";
        when 9927 => y_in <= "10100110"; x_in <= "01000111"; z_correct<="1110011100001010";
        when 9928 => y_in <= "10100110"; x_in <= "01001000"; z_correct<="1110011010110000";
        when 9929 => y_in <= "10100110"; x_in <= "01001001"; z_correct<="1110011001010110";
        when 9930 => y_in <= "10100110"; x_in <= "01001010"; z_correct<="1110010111111100";
        when 9931 => y_in <= "10100110"; x_in <= "01001011"; z_correct<="1110010110100010";
        when 9932 => y_in <= "10100110"; x_in <= "01001100"; z_correct<="1110010101001000";
        when 9933 => y_in <= "10100110"; x_in <= "01001101"; z_correct<="1110010011101110";
        when 9934 => y_in <= "10100110"; x_in <= "01001110"; z_correct<="1110010010010100";
        when 9935 => y_in <= "10100110"; x_in <= "01001111"; z_correct<="1110010000111010";
        when 9936 => y_in <= "10100110"; x_in <= "01010000"; z_correct<="1110001111100000";
        when 9937 => y_in <= "10100110"; x_in <= "01010001"; z_correct<="1110001110000110";
        when 9938 => y_in <= "10100110"; x_in <= "01010010"; z_correct<="1110001100101100";
        when 9939 => y_in <= "10100110"; x_in <= "01010011"; z_correct<="1110001011010010";
        when 9940 => y_in <= "10100110"; x_in <= "01010100"; z_correct<="1110001001111000";
        when 9941 => y_in <= "10100110"; x_in <= "01010101"; z_correct<="1110001000011110";
        when 9942 => y_in <= "10100110"; x_in <= "01010110"; z_correct<="1110000111000100";
        when 9943 => y_in <= "10100110"; x_in <= "01010111"; z_correct<="1110000101101010";
        when 9944 => y_in <= "10100110"; x_in <= "01011000"; z_correct<="1110000100010000";
        when 9945 => y_in <= "10100110"; x_in <= "01011001"; z_correct<="1110000010110110";
        when 9946 => y_in <= "10100110"; x_in <= "01011010"; z_correct<="1110000001011100";
        when 9947 => y_in <= "10100110"; x_in <= "01011011"; z_correct<="1110000000000010";
        when 9948 => y_in <= "10100110"; x_in <= "01011100"; z_correct<="1101111110101000";
        when 9949 => y_in <= "10100110"; x_in <= "01011101"; z_correct<="1101111101001110";
        when 9950 => y_in <= "10100110"; x_in <= "01011110"; z_correct<="1101111011110100";
        when 9951 => y_in <= "10100110"; x_in <= "01011111"; z_correct<="1101111010011010";
        when 9952 => y_in <= "10100110"; x_in <= "01100000"; z_correct<="1101111001000000";
        when 9953 => y_in <= "10100110"; x_in <= "01100001"; z_correct<="1101110111100110";
        when 9954 => y_in <= "10100110"; x_in <= "01100010"; z_correct<="1101110110001100";
        when 9955 => y_in <= "10100110"; x_in <= "01100011"; z_correct<="1101110100110010";
        when 9956 => y_in <= "10100110"; x_in <= "01100100"; z_correct<="1101110011011000";
        when 9957 => y_in <= "10100110"; x_in <= "01100101"; z_correct<="1101110001111110";
        when 9958 => y_in <= "10100110"; x_in <= "01100110"; z_correct<="1101110000100100";
        when 9959 => y_in <= "10100110"; x_in <= "01100111"; z_correct<="1101101111001010";
        when 9960 => y_in <= "10100110"; x_in <= "01101000"; z_correct<="1101101101110000";
        when 9961 => y_in <= "10100110"; x_in <= "01101001"; z_correct<="1101101100010110";
        when 9962 => y_in <= "10100110"; x_in <= "01101010"; z_correct<="1101101010111100";
        when 9963 => y_in <= "10100110"; x_in <= "01101011"; z_correct<="1101101001100010";
        when 9964 => y_in <= "10100110"; x_in <= "01101100"; z_correct<="1101101000001000";
        when 9965 => y_in <= "10100110"; x_in <= "01101101"; z_correct<="1101100110101110";
        when 9966 => y_in <= "10100110"; x_in <= "01101110"; z_correct<="1101100101010100";
        when 9967 => y_in <= "10100110"; x_in <= "01101111"; z_correct<="1101100011111010";
        when 9968 => y_in <= "10100110"; x_in <= "01110000"; z_correct<="1101100010100000";
        when 9969 => y_in <= "10100110"; x_in <= "01110001"; z_correct<="1101100001000110";
        when 9970 => y_in <= "10100110"; x_in <= "01110010"; z_correct<="1101011111101100";
        when 9971 => y_in <= "10100110"; x_in <= "01110011"; z_correct<="1101011110010010";
        when 9972 => y_in <= "10100110"; x_in <= "01110100"; z_correct<="1101011100111000";
        when 9973 => y_in <= "10100110"; x_in <= "01110101"; z_correct<="1101011011011110";
        when 9974 => y_in <= "10100110"; x_in <= "01110110"; z_correct<="1101011010000100";
        when 9975 => y_in <= "10100110"; x_in <= "01110111"; z_correct<="1101011000101010";
        when 9976 => y_in <= "10100110"; x_in <= "01111000"; z_correct<="1101010111010000";
        when 9977 => y_in <= "10100110"; x_in <= "01111001"; z_correct<="1101010101110110";
        when 9978 => y_in <= "10100110"; x_in <= "01111010"; z_correct<="1101010100011100";
        when 9979 => y_in <= "10100110"; x_in <= "01111011"; z_correct<="1101010011000010";
        when 9980 => y_in <= "10100110"; x_in <= "01111100"; z_correct<="1101010001101000";
        when 9981 => y_in <= "10100110"; x_in <= "01111101"; z_correct<="1101010000001110";
        when 9982 => y_in <= "10100110"; x_in <= "01111110"; z_correct<="1101001110110100";
        when 9983 => y_in <= "10100110"; x_in <= "01111111"; z_correct<="1101001101011010";
        when 9984 => y_in <= "10100111"; x_in <= "10000000"; z_correct<="0010110010000000";
        when 9985 => y_in <= "10100111"; x_in <= "10000001"; z_correct<="0010110000100111";
        when 9986 => y_in <= "10100111"; x_in <= "10000010"; z_correct<="0010101111001110";
        when 9987 => y_in <= "10100111"; x_in <= "10000011"; z_correct<="0010101101110101";
        when 9988 => y_in <= "10100111"; x_in <= "10000100"; z_correct<="0010101100011100";
        when 9989 => y_in <= "10100111"; x_in <= "10000101"; z_correct<="0010101011000011";
        when 9990 => y_in <= "10100111"; x_in <= "10000110"; z_correct<="0010101001101010";
        when 9991 => y_in <= "10100111"; x_in <= "10000111"; z_correct<="0010101000010001";
        when 9992 => y_in <= "10100111"; x_in <= "10001000"; z_correct<="0010100110111000";
        when 9993 => y_in <= "10100111"; x_in <= "10001001"; z_correct<="0010100101011111";
        when 9994 => y_in <= "10100111"; x_in <= "10001010"; z_correct<="0010100100000110";
        when 9995 => y_in <= "10100111"; x_in <= "10001011"; z_correct<="0010100010101101";
        when 9996 => y_in <= "10100111"; x_in <= "10001100"; z_correct<="0010100001010100";
        when 9997 => y_in <= "10100111"; x_in <= "10001101"; z_correct<="0010011111111011";
        when 9998 => y_in <= "10100111"; x_in <= "10001110"; z_correct<="0010011110100010";
        when 9999 => y_in <= "10100111"; x_in <= "10001111"; z_correct<="0010011101001001";
        when 10000 => y_in <= "10100111"; x_in <= "10010000"; z_correct<="0010011011110000";
        when 10001 => y_in <= "10100111"; x_in <= "10010001"; z_correct<="0010011010010111";
        when 10002 => y_in <= "10100111"; x_in <= "10010010"; z_correct<="0010011000111110";
        when 10003 => y_in <= "10100111"; x_in <= "10010011"; z_correct<="0010010111100101";
        when 10004 => y_in <= "10100111"; x_in <= "10010100"; z_correct<="0010010110001100";
        when 10005 => y_in <= "10100111"; x_in <= "10010101"; z_correct<="0010010100110011";
        when 10006 => y_in <= "10100111"; x_in <= "10010110"; z_correct<="0010010011011010";
        when 10007 => y_in <= "10100111"; x_in <= "10010111"; z_correct<="0010010010000001";
        when 10008 => y_in <= "10100111"; x_in <= "10011000"; z_correct<="0010010000101000";
        when 10009 => y_in <= "10100111"; x_in <= "10011001"; z_correct<="0010001111001111";
        when 10010 => y_in <= "10100111"; x_in <= "10011010"; z_correct<="0010001101110110";
        when 10011 => y_in <= "10100111"; x_in <= "10011011"; z_correct<="0010001100011101";
        when 10012 => y_in <= "10100111"; x_in <= "10011100"; z_correct<="0010001011000100";
        when 10013 => y_in <= "10100111"; x_in <= "10011101"; z_correct<="0010001001101011";
        when 10014 => y_in <= "10100111"; x_in <= "10011110"; z_correct<="0010001000010010";
        when 10015 => y_in <= "10100111"; x_in <= "10011111"; z_correct<="0010000110111001";
        when 10016 => y_in <= "10100111"; x_in <= "10100000"; z_correct<="0010000101100000";
        when 10017 => y_in <= "10100111"; x_in <= "10100001"; z_correct<="0010000100000111";
        when 10018 => y_in <= "10100111"; x_in <= "10100010"; z_correct<="0010000010101110";
        when 10019 => y_in <= "10100111"; x_in <= "10100011"; z_correct<="0010000001010101";
        when 10020 => y_in <= "10100111"; x_in <= "10100100"; z_correct<="0001111111111100";
        when 10021 => y_in <= "10100111"; x_in <= "10100101"; z_correct<="0001111110100011";
        when 10022 => y_in <= "10100111"; x_in <= "10100110"; z_correct<="0001111101001010";
        when 10023 => y_in <= "10100111"; x_in <= "10100111"; z_correct<="0001111011110001";
        when 10024 => y_in <= "10100111"; x_in <= "10101000"; z_correct<="0001111010011000";
        when 10025 => y_in <= "10100111"; x_in <= "10101001"; z_correct<="0001111000111111";
        when 10026 => y_in <= "10100111"; x_in <= "10101010"; z_correct<="0001110111100110";
        when 10027 => y_in <= "10100111"; x_in <= "10101011"; z_correct<="0001110110001101";
        when 10028 => y_in <= "10100111"; x_in <= "10101100"; z_correct<="0001110100110100";
        when 10029 => y_in <= "10100111"; x_in <= "10101101"; z_correct<="0001110011011011";
        when 10030 => y_in <= "10100111"; x_in <= "10101110"; z_correct<="0001110010000010";
        when 10031 => y_in <= "10100111"; x_in <= "10101111"; z_correct<="0001110000101001";
        when 10032 => y_in <= "10100111"; x_in <= "10110000"; z_correct<="0001101111010000";
        when 10033 => y_in <= "10100111"; x_in <= "10110001"; z_correct<="0001101101110111";
        when 10034 => y_in <= "10100111"; x_in <= "10110010"; z_correct<="0001101100011110";
        when 10035 => y_in <= "10100111"; x_in <= "10110011"; z_correct<="0001101011000101";
        when 10036 => y_in <= "10100111"; x_in <= "10110100"; z_correct<="0001101001101100";
        when 10037 => y_in <= "10100111"; x_in <= "10110101"; z_correct<="0001101000010011";
        when 10038 => y_in <= "10100111"; x_in <= "10110110"; z_correct<="0001100110111010";
        when 10039 => y_in <= "10100111"; x_in <= "10110111"; z_correct<="0001100101100001";
        when 10040 => y_in <= "10100111"; x_in <= "10111000"; z_correct<="0001100100001000";
        when 10041 => y_in <= "10100111"; x_in <= "10111001"; z_correct<="0001100010101111";
        when 10042 => y_in <= "10100111"; x_in <= "10111010"; z_correct<="0001100001010110";
        when 10043 => y_in <= "10100111"; x_in <= "10111011"; z_correct<="0001011111111101";
        when 10044 => y_in <= "10100111"; x_in <= "10111100"; z_correct<="0001011110100100";
        when 10045 => y_in <= "10100111"; x_in <= "10111101"; z_correct<="0001011101001011";
        when 10046 => y_in <= "10100111"; x_in <= "10111110"; z_correct<="0001011011110010";
        when 10047 => y_in <= "10100111"; x_in <= "10111111"; z_correct<="0001011010011001";
        when 10048 => y_in <= "10100111"; x_in <= "11000000"; z_correct<="0001011001000000";
        when 10049 => y_in <= "10100111"; x_in <= "11000001"; z_correct<="0001010111100111";
        when 10050 => y_in <= "10100111"; x_in <= "11000010"; z_correct<="0001010110001110";
        when 10051 => y_in <= "10100111"; x_in <= "11000011"; z_correct<="0001010100110101";
        when 10052 => y_in <= "10100111"; x_in <= "11000100"; z_correct<="0001010011011100";
        when 10053 => y_in <= "10100111"; x_in <= "11000101"; z_correct<="0001010010000011";
        when 10054 => y_in <= "10100111"; x_in <= "11000110"; z_correct<="0001010000101010";
        when 10055 => y_in <= "10100111"; x_in <= "11000111"; z_correct<="0001001111010001";
        when 10056 => y_in <= "10100111"; x_in <= "11001000"; z_correct<="0001001101111000";
        when 10057 => y_in <= "10100111"; x_in <= "11001001"; z_correct<="0001001100011111";
        when 10058 => y_in <= "10100111"; x_in <= "11001010"; z_correct<="0001001011000110";
        when 10059 => y_in <= "10100111"; x_in <= "11001011"; z_correct<="0001001001101101";
        when 10060 => y_in <= "10100111"; x_in <= "11001100"; z_correct<="0001001000010100";
        when 10061 => y_in <= "10100111"; x_in <= "11001101"; z_correct<="0001000110111011";
        when 10062 => y_in <= "10100111"; x_in <= "11001110"; z_correct<="0001000101100010";
        when 10063 => y_in <= "10100111"; x_in <= "11001111"; z_correct<="0001000100001001";
        when 10064 => y_in <= "10100111"; x_in <= "11010000"; z_correct<="0001000010110000";
        when 10065 => y_in <= "10100111"; x_in <= "11010001"; z_correct<="0001000001010111";
        when 10066 => y_in <= "10100111"; x_in <= "11010010"; z_correct<="0000111111111110";
        when 10067 => y_in <= "10100111"; x_in <= "11010011"; z_correct<="0000111110100101";
        when 10068 => y_in <= "10100111"; x_in <= "11010100"; z_correct<="0000111101001100";
        when 10069 => y_in <= "10100111"; x_in <= "11010101"; z_correct<="0000111011110011";
        when 10070 => y_in <= "10100111"; x_in <= "11010110"; z_correct<="0000111010011010";
        when 10071 => y_in <= "10100111"; x_in <= "11010111"; z_correct<="0000111001000001";
        when 10072 => y_in <= "10100111"; x_in <= "11011000"; z_correct<="0000110111101000";
        when 10073 => y_in <= "10100111"; x_in <= "11011001"; z_correct<="0000110110001111";
        when 10074 => y_in <= "10100111"; x_in <= "11011010"; z_correct<="0000110100110110";
        when 10075 => y_in <= "10100111"; x_in <= "11011011"; z_correct<="0000110011011101";
        when 10076 => y_in <= "10100111"; x_in <= "11011100"; z_correct<="0000110010000100";
        when 10077 => y_in <= "10100111"; x_in <= "11011101"; z_correct<="0000110000101011";
        when 10078 => y_in <= "10100111"; x_in <= "11011110"; z_correct<="0000101111010010";
        when 10079 => y_in <= "10100111"; x_in <= "11011111"; z_correct<="0000101101111001";
        when 10080 => y_in <= "10100111"; x_in <= "11100000"; z_correct<="0000101100100000";
        when 10081 => y_in <= "10100111"; x_in <= "11100001"; z_correct<="0000101011000111";
        when 10082 => y_in <= "10100111"; x_in <= "11100010"; z_correct<="0000101001101110";
        when 10083 => y_in <= "10100111"; x_in <= "11100011"; z_correct<="0000101000010101";
        when 10084 => y_in <= "10100111"; x_in <= "11100100"; z_correct<="0000100110111100";
        when 10085 => y_in <= "10100111"; x_in <= "11100101"; z_correct<="0000100101100011";
        when 10086 => y_in <= "10100111"; x_in <= "11100110"; z_correct<="0000100100001010";
        when 10087 => y_in <= "10100111"; x_in <= "11100111"; z_correct<="0000100010110001";
        when 10088 => y_in <= "10100111"; x_in <= "11101000"; z_correct<="0000100001011000";
        when 10089 => y_in <= "10100111"; x_in <= "11101001"; z_correct<="0000011111111111";
        when 10090 => y_in <= "10100111"; x_in <= "11101010"; z_correct<="0000011110100110";
        when 10091 => y_in <= "10100111"; x_in <= "11101011"; z_correct<="0000011101001101";
        when 10092 => y_in <= "10100111"; x_in <= "11101100"; z_correct<="0000011011110100";
        when 10093 => y_in <= "10100111"; x_in <= "11101101"; z_correct<="0000011010011011";
        when 10094 => y_in <= "10100111"; x_in <= "11101110"; z_correct<="0000011001000010";
        when 10095 => y_in <= "10100111"; x_in <= "11101111"; z_correct<="0000010111101001";
        when 10096 => y_in <= "10100111"; x_in <= "11110000"; z_correct<="0000010110010000";
        when 10097 => y_in <= "10100111"; x_in <= "11110001"; z_correct<="0000010100110111";
        when 10098 => y_in <= "10100111"; x_in <= "11110010"; z_correct<="0000010011011110";
        when 10099 => y_in <= "10100111"; x_in <= "11110011"; z_correct<="0000010010000101";
        when 10100 => y_in <= "10100111"; x_in <= "11110100"; z_correct<="0000010000101100";
        when 10101 => y_in <= "10100111"; x_in <= "11110101"; z_correct<="0000001111010011";
        when 10102 => y_in <= "10100111"; x_in <= "11110110"; z_correct<="0000001101111010";
        when 10103 => y_in <= "10100111"; x_in <= "11110111"; z_correct<="0000001100100001";
        when 10104 => y_in <= "10100111"; x_in <= "11111000"; z_correct<="0000001011001000";
        when 10105 => y_in <= "10100111"; x_in <= "11111001"; z_correct<="0000001001101111";
        when 10106 => y_in <= "10100111"; x_in <= "11111010"; z_correct<="0000001000010110";
        when 10107 => y_in <= "10100111"; x_in <= "11111011"; z_correct<="0000000110111101";
        when 10108 => y_in <= "10100111"; x_in <= "11111100"; z_correct<="0000000101100100";
        when 10109 => y_in <= "10100111"; x_in <= "11111101"; z_correct<="0000000100001011";
        when 10110 => y_in <= "10100111"; x_in <= "11111110"; z_correct<="0000000010110010";
        when 10111 => y_in <= "10100111"; x_in <= "11111111"; z_correct<="0000000001011001";
        when 10112 => y_in <= "10100111"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 10113 => y_in <= "10100111"; x_in <= "00000001"; z_correct<="1111111110100111";
        when 10114 => y_in <= "10100111"; x_in <= "00000010"; z_correct<="1111111101001110";
        when 10115 => y_in <= "10100111"; x_in <= "00000011"; z_correct<="1111111011110101";
        when 10116 => y_in <= "10100111"; x_in <= "00000100"; z_correct<="1111111010011100";
        when 10117 => y_in <= "10100111"; x_in <= "00000101"; z_correct<="1111111001000011";
        when 10118 => y_in <= "10100111"; x_in <= "00000110"; z_correct<="1111110111101010";
        when 10119 => y_in <= "10100111"; x_in <= "00000111"; z_correct<="1111110110010001";
        when 10120 => y_in <= "10100111"; x_in <= "00001000"; z_correct<="1111110100111000";
        when 10121 => y_in <= "10100111"; x_in <= "00001001"; z_correct<="1111110011011111";
        when 10122 => y_in <= "10100111"; x_in <= "00001010"; z_correct<="1111110010000110";
        when 10123 => y_in <= "10100111"; x_in <= "00001011"; z_correct<="1111110000101101";
        when 10124 => y_in <= "10100111"; x_in <= "00001100"; z_correct<="1111101111010100";
        when 10125 => y_in <= "10100111"; x_in <= "00001101"; z_correct<="1111101101111011";
        when 10126 => y_in <= "10100111"; x_in <= "00001110"; z_correct<="1111101100100010";
        when 10127 => y_in <= "10100111"; x_in <= "00001111"; z_correct<="1111101011001001";
        when 10128 => y_in <= "10100111"; x_in <= "00010000"; z_correct<="1111101001110000";
        when 10129 => y_in <= "10100111"; x_in <= "00010001"; z_correct<="1111101000010111";
        when 10130 => y_in <= "10100111"; x_in <= "00010010"; z_correct<="1111100110111110";
        when 10131 => y_in <= "10100111"; x_in <= "00010011"; z_correct<="1111100101100101";
        when 10132 => y_in <= "10100111"; x_in <= "00010100"; z_correct<="1111100100001100";
        when 10133 => y_in <= "10100111"; x_in <= "00010101"; z_correct<="1111100010110011";
        when 10134 => y_in <= "10100111"; x_in <= "00010110"; z_correct<="1111100001011010";
        when 10135 => y_in <= "10100111"; x_in <= "00010111"; z_correct<="1111100000000001";
        when 10136 => y_in <= "10100111"; x_in <= "00011000"; z_correct<="1111011110101000";
        when 10137 => y_in <= "10100111"; x_in <= "00011001"; z_correct<="1111011101001111";
        when 10138 => y_in <= "10100111"; x_in <= "00011010"; z_correct<="1111011011110110";
        when 10139 => y_in <= "10100111"; x_in <= "00011011"; z_correct<="1111011010011101";
        when 10140 => y_in <= "10100111"; x_in <= "00011100"; z_correct<="1111011001000100";
        when 10141 => y_in <= "10100111"; x_in <= "00011101"; z_correct<="1111010111101011";
        when 10142 => y_in <= "10100111"; x_in <= "00011110"; z_correct<="1111010110010010";
        when 10143 => y_in <= "10100111"; x_in <= "00011111"; z_correct<="1111010100111001";
        when 10144 => y_in <= "10100111"; x_in <= "00100000"; z_correct<="1111010011100000";
        when 10145 => y_in <= "10100111"; x_in <= "00100001"; z_correct<="1111010010000111";
        when 10146 => y_in <= "10100111"; x_in <= "00100010"; z_correct<="1111010000101110";
        when 10147 => y_in <= "10100111"; x_in <= "00100011"; z_correct<="1111001111010101";
        when 10148 => y_in <= "10100111"; x_in <= "00100100"; z_correct<="1111001101111100";
        when 10149 => y_in <= "10100111"; x_in <= "00100101"; z_correct<="1111001100100011";
        when 10150 => y_in <= "10100111"; x_in <= "00100110"; z_correct<="1111001011001010";
        when 10151 => y_in <= "10100111"; x_in <= "00100111"; z_correct<="1111001001110001";
        when 10152 => y_in <= "10100111"; x_in <= "00101000"; z_correct<="1111001000011000";
        when 10153 => y_in <= "10100111"; x_in <= "00101001"; z_correct<="1111000110111111";
        when 10154 => y_in <= "10100111"; x_in <= "00101010"; z_correct<="1111000101100110";
        when 10155 => y_in <= "10100111"; x_in <= "00101011"; z_correct<="1111000100001101";
        when 10156 => y_in <= "10100111"; x_in <= "00101100"; z_correct<="1111000010110100";
        when 10157 => y_in <= "10100111"; x_in <= "00101101"; z_correct<="1111000001011011";
        when 10158 => y_in <= "10100111"; x_in <= "00101110"; z_correct<="1111000000000010";
        when 10159 => y_in <= "10100111"; x_in <= "00101111"; z_correct<="1110111110101001";
        when 10160 => y_in <= "10100111"; x_in <= "00110000"; z_correct<="1110111101010000";
        when 10161 => y_in <= "10100111"; x_in <= "00110001"; z_correct<="1110111011110111";
        when 10162 => y_in <= "10100111"; x_in <= "00110010"; z_correct<="1110111010011110";
        when 10163 => y_in <= "10100111"; x_in <= "00110011"; z_correct<="1110111001000101";
        when 10164 => y_in <= "10100111"; x_in <= "00110100"; z_correct<="1110110111101100";
        when 10165 => y_in <= "10100111"; x_in <= "00110101"; z_correct<="1110110110010011";
        when 10166 => y_in <= "10100111"; x_in <= "00110110"; z_correct<="1110110100111010";
        when 10167 => y_in <= "10100111"; x_in <= "00110111"; z_correct<="1110110011100001";
        when 10168 => y_in <= "10100111"; x_in <= "00111000"; z_correct<="1110110010001000";
        when 10169 => y_in <= "10100111"; x_in <= "00111001"; z_correct<="1110110000101111";
        when 10170 => y_in <= "10100111"; x_in <= "00111010"; z_correct<="1110101111010110";
        when 10171 => y_in <= "10100111"; x_in <= "00111011"; z_correct<="1110101101111101";
        when 10172 => y_in <= "10100111"; x_in <= "00111100"; z_correct<="1110101100100100";
        when 10173 => y_in <= "10100111"; x_in <= "00111101"; z_correct<="1110101011001011";
        when 10174 => y_in <= "10100111"; x_in <= "00111110"; z_correct<="1110101001110010";
        when 10175 => y_in <= "10100111"; x_in <= "00111111"; z_correct<="1110101000011001";
        when 10176 => y_in <= "10100111"; x_in <= "01000000"; z_correct<="1110100111000000";
        when 10177 => y_in <= "10100111"; x_in <= "01000001"; z_correct<="1110100101100111";
        when 10178 => y_in <= "10100111"; x_in <= "01000010"; z_correct<="1110100100001110";
        when 10179 => y_in <= "10100111"; x_in <= "01000011"; z_correct<="1110100010110101";
        when 10180 => y_in <= "10100111"; x_in <= "01000100"; z_correct<="1110100001011100";
        when 10181 => y_in <= "10100111"; x_in <= "01000101"; z_correct<="1110100000000011";
        when 10182 => y_in <= "10100111"; x_in <= "01000110"; z_correct<="1110011110101010";
        when 10183 => y_in <= "10100111"; x_in <= "01000111"; z_correct<="1110011101010001";
        when 10184 => y_in <= "10100111"; x_in <= "01001000"; z_correct<="1110011011111000";
        when 10185 => y_in <= "10100111"; x_in <= "01001001"; z_correct<="1110011010011111";
        when 10186 => y_in <= "10100111"; x_in <= "01001010"; z_correct<="1110011001000110";
        when 10187 => y_in <= "10100111"; x_in <= "01001011"; z_correct<="1110010111101101";
        when 10188 => y_in <= "10100111"; x_in <= "01001100"; z_correct<="1110010110010100";
        when 10189 => y_in <= "10100111"; x_in <= "01001101"; z_correct<="1110010100111011";
        when 10190 => y_in <= "10100111"; x_in <= "01001110"; z_correct<="1110010011100010";
        when 10191 => y_in <= "10100111"; x_in <= "01001111"; z_correct<="1110010010001001";
        when 10192 => y_in <= "10100111"; x_in <= "01010000"; z_correct<="1110010000110000";
        when 10193 => y_in <= "10100111"; x_in <= "01010001"; z_correct<="1110001111010111";
        when 10194 => y_in <= "10100111"; x_in <= "01010010"; z_correct<="1110001101111110";
        when 10195 => y_in <= "10100111"; x_in <= "01010011"; z_correct<="1110001100100101";
        when 10196 => y_in <= "10100111"; x_in <= "01010100"; z_correct<="1110001011001100";
        when 10197 => y_in <= "10100111"; x_in <= "01010101"; z_correct<="1110001001110011";
        when 10198 => y_in <= "10100111"; x_in <= "01010110"; z_correct<="1110001000011010";
        when 10199 => y_in <= "10100111"; x_in <= "01010111"; z_correct<="1110000111000001";
        when 10200 => y_in <= "10100111"; x_in <= "01011000"; z_correct<="1110000101101000";
        when 10201 => y_in <= "10100111"; x_in <= "01011001"; z_correct<="1110000100001111";
        when 10202 => y_in <= "10100111"; x_in <= "01011010"; z_correct<="1110000010110110";
        when 10203 => y_in <= "10100111"; x_in <= "01011011"; z_correct<="1110000001011101";
        when 10204 => y_in <= "10100111"; x_in <= "01011100"; z_correct<="1110000000000100";
        when 10205 => y_in <= "10100111"; x_in <= "01011101"; z_correct<="1101111110101011";
        when 10206 => y_in <= "10100111"; x_in <= "01011110"; z_correct<="1101111101010010";
        when 10207 => y_in <= "10100111"; x_in <= "01011111"; z_correct<="1101111011111001";
        when 10208 => y_in <= "10100111"; x_in <= "01100000"; z_correct<="1101111010100000";
        when 10209 => y_in <= "10100111"; x_in <= "01100001"; z_correct<="1101111001000111";
        when 10210 => y_in <= "10100111"; x_in <= "01100010"; z_correct<="1101110111101110";
        when 10211 => y_in <= "10100111"; x_in <= "01100011"; z_correct<="1101110110010101";
        when 10212 => y_in <= "10100111"; x_in <= "01100100"; z_correct<="1101110100111100";
        when 10213 => y_in <= "10100111"; x_in <= "01100101"; z_correct<="1101110011100011";
        when 10214 => y_in <= "10100111"; x_in <= "01100110"; z_correct<="1101110010001010";
        when 10215 => y_in <= "10100111"; x_in <= "01100111"; z_correct<="1101110000110001";
        when 10216 => y_in <= "10100111"; x_in <= "01101000"; z_correct<="1101101111011000";
        when 10217 => y_in <= "10100111"; x_in <= "01101001"; z_correct<="1101101101111111";
        when 10218 => y_in <= "10100111"; x_in <= "01101010"; z_correct<="1101101100100110";
        when 10219 => y_in <= "10100111"; x_in <= "01101011"; z_correct<="1101101011001101";
        when 10220 => y_in <= "10100111"; x_in <= "01101100"; z_correct<="1101101001110100";
        when 10221 => y_in <= "10100111"; x_in <= "01101101"; z_correct<="1101101000011011";
        when 10222 => y_in <= "10100111"; x_in <= "01101110"; z_correct<="1101100111000010";
        when 10223 => y_in <= "10100111"; x_in <= "01101111"; z_correct<="1101100101101001";
        when 10224 => y_in <= "10100111"; x_in <= "01110000"; z_correct<="1101100100010000";
        when 10225 => y_in <= "10100111"; x_in <= "01110001"; z_correct<="1101100010110111";
        when 10226 => y_in <= "10100111"; x_in <= "01110010"; z_correct<="1101100001011110";
        when 10227 => y_in <= "10100111"; x_in <= "01110011"; z_correct<="1101100000000101";
        when 10228 => y_in <= "10100111"; x_in <= "01110100"; z_correct<="1101011110101100";
        when 10229 => y_in <= "10100111"; x_in <= "01110101"; z_correct<="1101011101010011";
        when 10230 => y_in <= "10100111"; x_in <= "01110110"; z_correct<="1101011011111010";
        when 10231 => y_in <= "10100111"; x_in <= "01110111"; z_correct<="1101011010100001";
        when 10232 => y_in <= "10100111"; x_in <= "01111000"; z_correct<="1101011001001000";
        when 10233 => y_in <= "10100111"; x_in <= "01111001"; z_correct<="1101010111101111";
        when 10234 => y_in <= "10100111"; x_in <= "01111010"; z_correct<="1101010110010110";
        when 10235 => y_in <= "10100111"; x_in <= "01111011"; z_correct<="1101010100111101";
        when 10236 => y_in <= "10100111"; x_in <= "01111100"; z_correct<="1101010011100100";
        when 10237 => y_in <= "10100111"; x_in <= "01111101"; z_correct<="1101010010001011";
        when 10238 => y_in <= "10100111"; x_in <= "01111110"; z_correct<="1101010000110010";
        when 10239 => y_in <= "10100111"; x_in <= "01111111"; z_correct<="1101001111011001";
        when 10240 => y_in <= "10101000"; x_in <= "10000000"; z_correct<="0010110000000000";
        when 10241 => y_in <= "10101000"; x_in <= "10000001"; z_correct<="0010101110101000";
        when 10242 => y_in <= "10101000"; x_in <= "10000010"; z_correct<="0010101101010000";
        when 10243 => y_in <= "10101000"; x_in <= "10000011"; z_correct<="0010101011111000";
        when 10244 => y_in <= "10101000"; x_in <= "10000100"; z_correct<="0010101010100000";
        when 10245 => y_in <= "10101000"; x_in <= "10000101"; z_correct<="0010101001001000";
        when 10246 => y_in <= "10101000"; x_in <= "10000110"; z_correct<="0010100111110000";
        when 10247 => y_in <= "10101000"; x_in <= "10000111"; z_correct<="0010100110011000";
        when 10248 => y_in <= "10101000"; x_in <= "10001000"; z_correct<="0010100101000000";
        when 10249 => y_in <= "10101000"; x_in <= "10001001"; z_correct<="0010100011101000";
        when 10250 => y_in <= "10101000"; x_in <= "10001010"; z_correct<="0010100010010000";
        when 10251 => y_in <= "10101000"; x_in <= "10001011"; z_correct<="0010100000111000";
        when 10252 => y_in <= "10101000"; x_in <= "10001100"; z_correct<="0010011111100000";
        when 10253 => y_in <= "10101000"; x_in <= "10001101"; z_correct<="0010011110001000";
        when 10254 => y_in <= "10101000"; x_in <= "10001110"; z_correct<="0010011100110000";
        when 10255 => y_in <= "10101000"; x_in <= "10001111"; z_correct<="0010011011011000";
        when 10256 => y_in <= "10101000"; x_in <= "10010000"; z_correct<="0010011010000000";
        when 10257 => y_in <= "10101000"; x_in <= "10010001"; z_correct<="0010011000101000";
        when 10258 => y_in <= "10101000"; x_in <= "10010010"; z_correct<="0010010111010000";
        when 10259 => y_in <= "10101000"; x_in <= "10010011"; z_correct<="0010010101111000";
        when 10260 => y_in <= "10101000"; x_in <= "10010100"; z_correct<="0010010100100000";
        when 10261 => y_in <= "10101000"; x_in <= "10010101"; z_correct<="0010010011001000";
        when 10262 => y_in <= "10101000"; x_in <= "10010110"; z_correct<="0010010001110000";
        when 10263 => y_in <= "10101000"; x_in <= "10010111"; z_correct<="0010010000011000";
        when 10264 => y_in <= "10101000"; x_in <= "10011000"; z_correct<="0010001111000000";
        when 10265 => y_in <= "10101000"; x_in <= "10011001"; z_correct<="0010001101101000";
        when 10266 => y_in <= "10101000"; x_in <= "10011010"; z_correct<="0010001100010000";
        when 10267 => y_in <= "10101000"; x_in <= "10011011"; z_correct<="0010001010111000";
        when 10268 => y_in <= "10101000"; x_in <= "10011100"; z_correct<="0010001001100000";
        when 10269 => y_in <= "10101000"; x_in <= "10011101"; z_correct<="0010001000001000";
        when 10270 => y_in <= "10101000"; x_in <= "10011110"; z_correct<="0010000110110000";
        when 10271 => y_in <= "10101000"; x_in <= "10011111"; z_correct<="0010000101011000";
        when 10272 => y_in <= "10101000"; x_in <= "10100000"; z_correct<="0010000100000000";
        when 10273 => y_in <= "10101000"; x_in <= "10100001"; z_correct<="0010000010101000";
        when 10274 => y_in <= "10101000"; x_in <= "10100010"; z_correct<="0010000001010000";
        when 10275 => y_in <= "10101000"; x_in <= "10100011"; z_correct<="0001111111111000";
        when 10276 => y_in <= "10101000"; x_in <= "10100100"; z_correct<="0001111110100000";
        when 10277 => y_in <= "10101000"; x_in <= "10100101"; z_correct<="0001111101001000";
        when 10278 => y_in <= "10101000"; x_in <= "10100110"; z_correct<="0001111011110000";
        when 10279 => y_in <= "10101000"; x_in <= "10100111"; z_correct<="0001111010011000";
        when 10280 => y_in <= "10101000"; x_in <= "10101000"; z_correct<="0001111001000000";
        when 10281 => y_in <= "10101000"; x_in <= "10101001"; z_correct<="0001110111101000";
        when 10282 => y_in <= "10101000"; x_in <= "10101010"; z_correct<="0001110110010000";
        when 10283 => y_in <= "10101000"; x_in <= "10101011"; z_correct<="0001110100111000";
        when 10284 => y_in <= "10101000"; x_in <= "10101100"; z_correct<="0001110011100000";
        when 10285 => y_in <= "10101000"; x_in <= "10101101"; z_correct<="0001110010001000";
        when 10286 => y_in <= "10101000"; x_in <= "10101110"; z_correct<="0001110000110000";
        when 10287 => y_in <= "10101000"; x_in <= "10101111"; z_correct<="0001101111011000";
        when 10288 => y_in <= "10101000"; x_in <= "10110000"; z_correct<="0001101110000000";
        when 10289 => y_in <= "10101000"; x_in <= "10110001"; z_correct<="0001101100101000";
        when 10290 => y_in <= "10101000"; x_in <= "10110010"; z_correct<="0001101011010000";
        when 10291 => y_in <= "10101000"; x_in <= "10110011"; z_correct<="0001101001111000";
        when 10292 => y_in <= "10101000"; x_in <= "10110100"; z_correct<="0001101000100000";
        when 10293 => y_in <= "10101000"; x_in <= "10110101"; z_correct<="0001100111001000";
        when 10294 => y_in <= "10101000"; x_in <= "10110110"; z_correct<="0001100101110000";
        when 10295 => y_in <= "10101000"; x_in <= "10110111"; z_correct<="0001100100011000";
        when 10296 => y_in <= "10101000"; x_in <= "10111000"; z_correct<="0001100011000000";
        when 10297 => y_in <= "10101000"; x_in <= "10111001"; z_correct<="0001100001101000";
        when 10298 => y_in <= "10101000"; x_in <= "10111010"; z_correct<="0001100000010000";
        when 10299 => y_in <= "10101000"; x_in <= "10111011"; z_correct<="0001011110111000";
        when 10300 => y_in <= "10101000"; x_in <= "10111100"; z_correct<="0001011101100000";
        when 10301 => y_in <= "10101000"; x_in <= "10111101"; z_correct<="0001011100001000";
        when 10302 => y_in <= "10101000"; x_in <= "10111110"; z_correct<="0001011010110000";
        when 10303 => y_in <= "10101000"; x_in <= "10111111"; z_correct<="0001011001011000";
        when 10304 => y_in <= "10101000"; x_in <= "11000000"; z_correct<="0001011000000000";
        when 10305 => y_in <= "10101000"; x_in <= "11000001"; z_correct<="0001010110101000";
        when 10306 => y_in <= "10101000"; x_in <= "11000010"; z_correct<="0001010101010000";
        when 10307 => y_in <= "10101000"; x_in <= "11000011"; z_correct<="0001010011111000";
        when 10308 => y_in <= "10101000"; x_in <= "11000100"; z_correct<="0001010010100000";
        when 10309 => y_in <= "10101000"; x_in <= "11000101"; z_correct<="0001010001001000";
        when 10310 => y_in <= "10101000"; x_in <= "11000110"; z_correct<="0001001111110000";
        when 10311 => y_in <= "10101000"; x_in <= "11000111"; z_correct<="0001001110011000";
        when 10312 => y_in <= "10101000"; x_in <= "11001000"; z_correct<="0001001101000000";
        when 10313 => y_in <= "10101000"; x_in <= "11001001"; z_correct<="0001001011101000";
        when 10314 => y_in <= "10101000"; x_in <= "11001010"; z_correct<="0001001010010000";
        when 10315 => y_in <= "10101000"; x_in <= "11001011"; z_correct<="0001001000111000";
        when 10316 => y_in <= "10101000"; x_in <= "11001100"; z_correct<="0001000111100000";
        when 10317 => y_in <= "10101000"; x_in <= "11001101"; z_correct<="0001000110001000";
        when 10318 => y_in <= "10101000"; x_in <= "11001110"; z_correct<="0001000100110000";
        when 10319 => y_in <= "10101000"; x_in <= "11001111"; z_correct<="0001000011011000";
        when 10320 => y_in <= "10101000"; x_in <= "11010000"; z_correct<="0001000010000000";
        when 10321 => y_in <= "10101000"; x_in <= "11010001"; z_correct<="0001000000101000";
        when 10322 => y_in <= "10101000"; x_in <= "11010010"; z_correct<="0000111111010000";
        when 10323 => y_in <= "10101000"; x_in <= "11010011"; z_correct<="0000111101111000";
        when 10324 => y_in <= "10101000"; x_in <= "11010100"; z_correct<="0000111100100000";
        when 10325 => y_in <= "10101000"; x_in <= "11010101"; z_correct<="0000111011001000";
        when 10326 => y_in <= "10101000"; x_in <= "11010110"; z_correct<="0000111001110000";
        when 10327 => y_in <= "10101000"; x_in <= "11010111"; z_correct<="0000111000011000";
        when 10328 => y_in <= "10101000"; x_in <= "11011000"; z_correct<="0000110111000000";
        when 10329 => y_in <= "10101000"; x_in <= "11011001"; z_correct<="0000110101101000";
        when 10330 => y_in <= "10101000"; x_in <= "11011010"; z_correct<="0000110100010000";
        when 10331 => y_in <= "10101000"; x_in <= "11011011"; z_correct<="0000110010111000";
        when 10332 => y_in <= "10101000"; x_in <= "11011100"; z_correct<="0000110001100000";
        when 10333 => y_in <= "10101000"; x_in <= "11011101"; z_correct<="0000110000001000";
        when 10334 => y_in <= "10101000"; x_in <= "11011110"; z_correct<="0000101110110000";
        when 10335 => y_in <= "10101000"; x_in <= "11011111"; z_correct<="0000101101011000";
        when 10336 => y_in <= "10101000"; x_in <= "11100000"; z_correct<="0000101100000000";
        when 10337 => y_in <= "10101000"; x_in <= "11100001"; z_correct<="0000101010101000";
        when 10338 => y_in <= "10101000"; x_in <= "11100010"; z_correct<="0000101001010000";
        when 10339 => y_in <= "10101000"; x_in <= "11100011"; z_correct<="0000100111111000";
        when 10340 => y_in <= "10101000"; x_in <= "11100100"; z_correct<="0000100110100000";
        when 10341 => y_in <= "10101000"; x_in <= "11100101"; z_correct<="0000100101001000";
        when 10342 => y_in <= "10101000"; x_in <= "11100110"; z_correct<="0000100011110000";
        when 10343 => y_in <= "10101000"; x_in <= "11100111"; z_correct<="0000100010011000";
        when 10344 => y_in <= "10101000"; x_in <= "11101000"; z_correct<="0000100001000000";
        when 10345 => y_in <= "10101000"; x_in <= "11101001"; z_correct<="0000011111101000";
        when 10346 => y_in <= "10101000"; x_in <= "11101010"; z_correct<="0000011110010000";
        when 10347 => y_in <= "10101000"; x_in <= "11101011"; z_correct<="0000011100111000";
        when 10348 => y_in <= "10101000"; x_in <= "11101100"; z_correct<="0000011011100000";
        when 10349 => y_in <= "10101000"; x_in <= "11101101"; z_correct<="0000011010001000";
        when 10350 => y_in <= "10101000"; x_in <= "11101110"; z_correct<="0000011000110000";
        when 10351 => y_in <= "10101000"; x_in <= "11101111"; z_correct<="0000010111011000";
        when 10352 => y_in <= "10101000"; x_in <= "11110000"; z_correct<="0000010110000000";
        when 10353 => y_in <= "10101000"; x_in <= "11110001"; z_correct<="0000010100101000";
        when 10354 => y_in <= "10101000"; x_in <= "11110010"; z_correct<="0000010011010000";
        when 10355 => y_in <= "10101000"; x_in <= "11110011"; z_correct<="0000010001111000";
        when 10356 => y_in <= "10101000"; x_in <= "11110100"; z_correct<="0000010000100000";
        when 10357 => y_in <= "10101000"; x_in <= "11110101"; z_correct<="0000001111001000";
        when 10358 => y_in <= "10101000"; x_in <= "11110110"; z_correct<="0000001101110000";
        when 10359 => y_in <= "10101000"; x_in <= "11110111"; z_correct<="0000001100011000";
        when 10360 => y_in <= "10101000"; x_in <= "11111000"; z_correct<="0000001011000000";
        when 10361 => y_in <= "10101000"; x_in <= "11111001"; z_correct<="0000001001101000";
        when 10362 => y_in <= "10101000"; x_in <= "11111010"; z_correct<="0000001000010000";
        when 10363 => y_in <= "10101000"; x_in <= "11111011"; z_correct<="0000000110111000";
        when 10364 => y_in <= "10101000"; x_in <= "11111100"; z_correct<="0000000101100000";
        when 10365 => y_in <= "10101000"; x_in <= "11111101"; z_correct<="0000000100001000";
        when 10366 => y_in <= "10101000"; x_in <= "11111110"; z_correct<="0000000010110000";
        when 10367 => y_in <= "10101000"; x_in <= "11111111"; z_correct<="0000000001011000";
        when 10368 => y_in <= "10101000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 10369 => y_in <= "10101000"; x_in <= "00000001"; z_correct<="1111111110101000";
        when 10370 => y_in <= "10101000"; x_in <= "00000010"; z_correct<="1111111101010000";
        when 10371 => y_in <= "10101000"; x_in <= "00000011"; z_correct<="1111111011111000";
        when 10372 => y_in <= "10101000"; x_in <= "00000100"; z_correct<="1111111010100000";
        when 10373 => y_in <= "10101000"; x_in <= "00000101"; z_correct<="1111111001001000";
        when 10374 => y_in <= "10101000"; x_in <= "00000110"; z_correct<="1111110111110000";
        when 10375 => y_in <= "10101000"; x_in <= "00000111"; z_correct<="1111110110011000";
        when 10376 => y_in <= "10101000"; x_in <= "00001000"; z_correct<="1111110101000000";
        when 10377 => y_in <= "10101000"; x_in <= "00001001"; z_correct<="1111110011101000";
        when 10378 => y_in <= "10101000"; x_in <= "00001010"; z_correct<="1111110010010000";
        when 10379 => y_in <= "10101000"; x_in <= "00001011"; z_correct<="1111110000111000";
        when 10380 => y_in <= "10101000"; x_in <= "00001100"; z_correct<="1111101111100000";
        when 10381 => y_in <= "10101000"; x_in <= "00001101"; z_correct<="1111101110001000";
        when 10382 => y_in <= "10101000"; x_in <= "00001110"; z_correct<="1111101100110000";
        when 10383 => y_in <= "10101000"; x_in <= "00001111"; z_correct<="1111101011011000";
        when 10384 => y_in <= "10101000"; x_in <= "00010000"; z_correct<="1111101010000000";
        when 10385 => y_in <= "10101000"; x_in <= "00010001"; z_correct<="1111101000101000";
        when 10386 => y_in <= "10101000"; x_in <= "00010010"; z_correct<="1111100111010000";
        when 10387 => y_in <= "10101000"; x_in <= "00010011"; z_correct<="1111100101111000";
        when 10388 => y_in <= "10101000"; x_in <= "00010100"; z_correct<="1111100100100000";
        when 10389 => y_in <= "10101000"; x_in <= "00010101"; z_correct<="1111100011001000";
        when 10390 => y_in <= "10101000"; x_in <= "00010110"; z_correct<="1111100001110000";
        when 10391 => y_in <= "10101000"; x_in <= "00010111"; z_correct<="1111100000011000";
        when 10392 => y_in <= "10101000"; x_in <= "00011000"; z_correct<="1111011111000000";
        when 10393 => y_in <= "10101000"; x_in <= "00011001"; z_correct<="1111011101101000";
        when 10394 => y_in <= "10101000"; x_in <= "00011010"; z_correct<="1111011100010000";
        when 10395 => y_in <= "10101000"; x_in <= "00011011"; z_correct<="1111011010111000";
        when 10396 => y_in <= "10101000"; x_in <= "00011100"; z_correct<="1111011001100000";
        when 10397 => y_in <= "10101000"; x_in <= "00011101"; z_correct<="1111011000001000";
        when 10398 => y_in <= "10101000"; x_in <= "00011110"; z_correct<="1111010110110000";
        when 10399 => y_in <= "10101000"; x_in <= "00011111"; z_correct<="1111010101011000";
        when 10400 => y_in <= "10101000"; x_in <= "00100000"; z_correct<="1111010100000000";
        when 10401 => y_in <= "10101000"; x_in <= "00100001"; z_correct<="1111010010101000";
        when 10402 => y_in <= "10101000"; x_in <= "00100010"; z_correct<="1111010001010000";
        when 10403 => y_in <= "10101000"; x_in <= "00100011"; z_correct<="1111001111111000";
        when 10404 => y_in <= "10101000"; x_in <= "00100100"; z_correct<="1111001110100000";
        when 10405 => y_in <= "10101000"; x_in <= "00100101"; z_correct<="1111001101001000";
        when 10406 => y_in <= "10101000"; x_in <= "00100110"; z_correct<="1111001011110000";
        when 10407 => y_in <= "10101000"; x_in <= "00100111"; z_correct<="1111001010011000";
        when 10408 => y_in <= "10101000"; x_in <= "00101000"; z_correct<="1111001001000000";
        when 10409 => y_in <= "10101000"; x_in <= "00101001"; z_correct<="1111000111101000";
        when 10410 => y_in <= "10101000"; x_in <= "00101010"; z_correct<="1111000110010000";
        when 10411 => y_in <= "10101000"; x_in <= "00101011"; z_correct<="1111000100111000";
        when 10412 => y_in <= "10101000"; x_in <= "00101100"; z_correct<="1111000011100000";
        when 10413 => y_in <= "10101000"; x_in <= "00101101"; z_correct<="1111000010001000";
        when 10414 => y_in <= "10101000"; x_in <= "00101110"; z_correct<="1111000000110000";
        when 10415 => y_in <= "10101000"; x_in <= "00101111"; z_correct<="1110111111011000";
        when 10416 => y_in <= "10101000"; x_in <= "00110000"; z_correct<="1110111110000000";
        when 10417 => y_in <= "10101000"; x_in <= "00110001"; z_correct<="1110111100101000";
        when 10418 => y_in <= "10101000"; x_in <= "00110010"; z_correct<="1110111011010000";
        when 10419 => y_in <= "10101000"; x_in <= "00110011"; z_correct<="1110111001111000";
        when 10420 => y_in <= "10101000"; x_in <= "00110100"; z_correct<="1110111000100000";
        when 10421 => y_in <= "10101000"; x_in <= "00110101"; z_correct<="1110110111001000";
        when 10422 => y_in <= "10101000"; x_in <= "00110110"; z_correct<="1110110101110000";
        when 10423 => y_in <= "10101000"; x_in <= "00110111"; z_correct<="1110110100011000";
        when 10424 => y_in <= "10101000"; x_in <= "00111000"; z_correct<="1110110011000000";
        when 10425 => y_in <= "10101000"; x_in <= "00111001"; z_correct<="1110110001101000";
        when 10426 => y_in <= "10101000"; x_in <= "00111010"; z_correct<="1110110000010000";
        when 10427 => y_in <= "10101000"; x_in <= "00111011"; z_correct<="1110101110111000";
        when 10428 => y_in <= "10101000"; x_in <= "00111100"; z_correct<="1110101101100000";
        when 10429 => y_in <= "10101000"; x_in <= "00111101"; z_correct<="1110101100001000";
        when 10430 => y_in <= "10101000"; x_in <= "00111110"; z_correct<="1110101010110000";
        when 10431 => y_in <= "10101000"; x_in <= "00111111"; z_correct<="1110101001011000";
        when 10432 => y_in <= "10101000"; x_in <= "01000000"; z_correct<="1110101000000000";
        when 10433 => y_in <= "10101000"; x_in <= "01000001"; z_correct<="1110100110101000";
        when 10434 => y_in <= "10101000"; x_in <= "01000010"; z_correct<="1110100101010000";
        when 10435 => y_in <= "10101000"; x_in <= "01000011"; z_correct<="1110100011111000";
        when 10436 => y_in <= "10101000"; x_in <= "01000100"; z_correct<="1110100010100000";
        when 10437 => y_in <= "10101000"; x_in <= "01000101"; z_correct<="1110100001001000";
        when 10438 => y_in <= "10101000"; x_in <= "01000110"; z_correct<="1110011111110000";
        when 10439 => y_in <= "10101000"; x_in <= "01000111"; z_correct<="1110011110011000";
        when 10440 => y_in <= "10101000"; x_in <= "01001000"; z_correct<="1110011101000000";
        when 10441 => y_in <= "10101000"; x_in <= "01001001"; z_correct<="1110011011101000";
        when 10442 => y_in <= "10101000"; x_in <= "01001010"; z_correct<="1110011010010000";
        when 10443 => y_in <= "10101000"; x_in <= "01001011"; z_correct<="1110011000111000";
        when 10444 => y_in <= "10101000"; x_in <= "01001100"; z_correct<="1110010111100000";
        when 10445 => y_in <= "10101000"; x_in <= "01001101"; z_correct<="1110010110001000";
        when 10446 => y_in <= "10101000"; x_in <= "01001110"; z_correct<="1110010100110000";
        when 10447 => y_in <= "10101000"; x_in <= "01001111"; z_correct<="1110010011011000";
        when 10448 => y_in <= "10101000"; x_in <= "01010000"; z_correct<="1110010010000000";
        when 10449 => y_in <= "10101000"; x_in <= "01010001"; z_correct<="1110010000101000";
        when 10450 => y_in <= "10101000"; x_in <= "01010010"; z_correct<="1110001111010000";
        when 10451 => y_in <= "10101000"; x_in <= "01010011"; z_correct<="1110001101111000";
        when 10452 => y_in <= "10101000"; x_in <= "01010100"; z_correct<="1110001100100000";
        when 10453 => y_in <= "10101000"; x_in <= "01010101"; z_correct<="1110001011001000";
        when 10454 => y_in <= "10101000"; x_in <= "01010110"; z_correct<="1110001001110000";
        when 10455 => y_in <= "10101000"; x_in <= "01010111"; z_correct<="1110001000011000";
        when 10456 => y_in <= "10101000"; x_in <= "01011000"; z_correct<="1110000111000000";
        when 10457 => y_in <= "10101000"; x_in <= "01011001"; z_correct<="1110000101101000";
        when 10458 => y_in <= "10101000"; x_in <= "01011010"; z_correct<="1110000100010000";
        when 10459 => y_in <= "10101000"; x_in <= "01011011"; z_correct<="1110000010111000";
        when 10460 => y_in <= "10101000"; x_in <= "01011100"; z_correct<="1110000001100000";
        when 10461 => y_in <= "10101000"; x_in <= "01011101"; z_correct<="1110000000001000";
        when 10462 => y_in <= "10101000"; x_in <= "01011110"; z_correct<="1101111110110000";
        when 10463 => y_in <= "10101000"; x_in <= "01011111"; z_correct<="1101111101011000";
        when 10464 => y_in <= "10101000"; x_in <= "01100000"; z_correct<="1101111100000000";
        when 10465 => y_in <= "10101000"; x_in <= "01100001"; z_correct<="1101111010101000";
        when 10466 => y_in <= "10101000"; x_in <= "01100010"; z_correct<="1101111001010000";
        when 10467 => y_in <= "10101000"; x_in <= "01100011"; z_correct<="1101110111111000";
        when 10468 => y_in <= "10101000"; x_in <= "01100100"; z_correct<="1101110110100000";
        when 10469 => y_in <= "10101000"; x_in <= "01100101"; z_correct<="1101110101001000";
        when 10470 => y_in <= "10101000"; x_in <= "01100110"; z_correct<="1101110011110000";
        when 10471 => y_in <= "10101000"; x_in <= "01100111"; z_correct<="1101110010011000";
        when 10472 => y_in <= "10101000"; x_in <= "01101000"; z_correct<="1101110001000000";
        when 10473 => y_in <= "10101000"; x_in <= "01101001"; z_correct<="1101101111101000";
        when 10474 => y_in <= "10101000"; x_in <= "01101010"; z_correct<="1101101110010000";
        when 10475 => y_in <= "10101000"; x_in <= "01101011"; z_correct<="1101101100111000";
        when 10476 => y_in <= "10101000"; x_in <= "01101100"; z_correct<="1101101011100000";
        when 10477 => y_in <= "10101000"; x_in <= "01101101"; z_correct<="1101101010001000";
        when 10478 => y_in <= "10101000"; x_in <= "01101110"; z_correct<="1101101000110000";
        when 10479 => y_in <= "10101000"; x_in <= "01101111"; z_correct<="1101100111011000";
        when 10480 => y_in <= "10101000"; x_in <= "01110000"; z_correct<="1101100110000000";
        when 10481 => y_in <= "10101000"; x_in <= "01110001"; z_correct<="1101100100101000";
        when 10482 => y_in <= "10101000"; x_in <= "01110010"; z_correct<="1101100011010000";
        when 10483 => y_in <= "10101000"; x_in <= "01110011"; z_correct<="1101100001111000";
        when 10484 => y_in <= "10101000"; x_in <= "01110100"; z_correct<="1101100000100000";
        when 10485 => y_in <= "10101000"; x_in <= "01110101"; z_correct<="1101011111001000";
        when 10486 => y_in <= "10101000"; x_in <= "01110110"; z_correct<="1101011101110000";
        when 10487 => y_in <= "10101000"; x_in <= "01110111"; z_correct<="1101011100011000";
        when 10488 => y_in <= "10101000"; x_in <= "01111000"; z_correct<="1101011011000000";
        when 10489 => y_in <= "10101000"; x_in <= "01111001"; z_correct<="1101011001101000";
        when 10490 => y_in <= "10101000"; x_in <= "01111010"; z_correct<="1101011000010000";
        when 10491 => y_in <= "10101000"; x_in <= "01111011"; z_correct<="1101010110111000";
        when 10492 => y_in <= "10101000"; x_in <= "01111100"; z_correct<="1101010101100000";
        when 10493 => y_in <= "10101000"; x_in <= "01111101"; z_correct<="1101010100001000";
        when 10494 => y_in <= "10101000"; x_in <= "01111110"; z_correct<="1101010010110000";
        when 10495 => y_in <= "10101000"; x_in <= "01111111"; z_correct<="1101010001011000";
        when 10496 => y_in <= "10101001"; x_in <= "10000000"; z_correct<="0010101110000000";
        when 10497 => y_in <= "10101001"; x_in <= "10000001"; z_correct<="0010101100101001";
        when 10498 => y_in <= "10101001"; x_in <= "10000010"; z_correct<="0010101011010010";
        when 10499 => y_in <= "10101001"; x_in <= "10000011"; z_correct<="0010101001111011";
        when 10500 => y_in <= "10101001"; x_in <= "10000100"; z_correct<="0010101000100100";
        when 10501 => y_in <= "10101001"; x_in <= "10000101"; z_correct<="0010100111001101";
        when 10502 => y_in <= "10101001"; x_in <= "10000110"; z_correct<="0010100101110110";
        when 10503 => y_in <= "10101001"; x_in <= "10000111"; z_correct<="0010100100011111";
        when 10504 => y_in <= "10101001"; x_in <= "10001000"; z_correct<="0010100011001000";
        when 10505 => y_in <= "10101001"; x_in <= "10001001"; z_correct<="0010100001110001";
        when 10506 => y_in <= "10101001"; x_in <= "10001010"; z_correct<="0010100000011010";
        when 10507 => y_in <= "10101001"; x_in <= "10001011"; z_correct<="0010011111000011";
        when 10508 => y_in <= "10101001"; x_in <= "10001100"; z_correct<="0010011101101100";
        when 10509 => y_in <= "10101001"; x_in <= "10001101"; z_correct<="0010011100010101";
        when 10510 => y_in <= "10101001"; x_in <= "10001110"; z_correct<="0010011010111110";
        when 10511 => y_in <= "10101001"; x_in <= "10001111"; z_correct<="0010011001100111";
        when 10512 => y_in <= "10101001"; x_in <= "10010000"; z_correct<="0010011000010000";
        when 10513 => y_in <= "10101001"; x_in <= "10010001"; z_correct<="0010010110111001";
        when 10514 => y_in <= "10101001"; x_in <= "10010010"; z_correct<="0010010101100010";
        when 10515 => y_in <= "10101001"; x_in <= "10010011"; z_correct<="0010010100001011";
        when 10516 => y_in <= "10101001"; x_in <= "10010100"; z_correct<="0010010010110100";
        when 10517 => y_in <= "10101001"; x_in <= "10010101"; z_correct<="0010010001011101";
        when 10518 => y_in <= "10101001"; x_in <= "10010110"; z_correct<="0010010000000110";
        when 10519 => y_in <= "10101001"; x_in <= "10010111"; z_correct<="0010001110101111";
        when 10520 => y_in <= "10101001"; x_in <= "10011000"; z_correct<="0010001101011000";
        when 10521 => y_in <= "10101001"; x_in <= "10011001"; z_correct<="0010001100000001";
        when 10522 => y_in <= "10101001"; x_in <= "10011010"; z_correct<="0010001010101010";
        when 10523 => y_in <= "10101001"; x_in <= "10011011"; z_correct<="0010001001010011";
        when 10524 => y_in <= "10101001"; x_in <= "10011100"; z_correct<="0010000111111100";
        when 10525 => y_in <= "10101001"; x_in <= "10011101"; z_correct<="0010000110100101";
        when 10526 => y_in <= "10101001"; x_in <= "10011110"; z_correct<="0010000101001110";
        when 10527 => y_in <= "10101001"; x_in <= "10011111"; z_correct<="0010000011110111";
        when 10528 => y_in <= "10101001"; x_in <= "10100000"; z_correct<="0010000010100000";
        when 10529 => y_in <= "10101001"; x_in <= "10100001"; z_correct<="0010000001001001";
        when 10530 => y_in <= "10101001"; x_in <= "10100010"; z_correct<="0001111111110010";
        when 10531 => y_in <= "10101001"; x_in <= "10100011"; z_correct<="0001111110011011";
        when 10532 => y_in <= "10101001"; x_in <= "10100100"; z_correct<="0001111101000100";
        when 10533 => y_in <= "10101001"; x_in <= "10100101"; z_correct<="0001111011101101";
        when 10534 => y_in <= "10101001"; x_in <= "10100110"; z_correct<="0001111010010110";
        when 10535 => y_in <= "10101001"; x_in <= "10100111"; z_correct<="0001111000111111";
        when 10536 => y_in <= "10101001"; x_in <= "10101000"; z_correct<="0001110111101000";
        when 10537 => y_in <= "10101001"; x_in <= "10101001"; z_correct<="0001110110010001";
        when 10538 => y_in <= "10101001"; x_in <= "10101010"; z_correct<="0001110100111010";
        when 10539 => y_in <= "10101001"; x_in <= "10101011"; z_correct<="0001110011100011";
        when 10540 => y_in <= "10101001"; x_in <= "10101100"; z_correct<="0001110010001100";
        when 10541 => y_in <= "10101001"; x_in <= "10101101"; z_correct<="0001110000110101";
        when 10542 => y_in <= "10101001"; x_in <= "10101110"; z_correct<="0001101111011110";
        when 10543 => y_in <= "10101001"; x_in <= "10101111"; z_correct<="0001101110000111";
        when 10544 => y_in <= "10101001"; x_in <= "10110000"; z_correct<="0001101100110000";
        when 10545 => y_in <= "10101001"; x_in <= "10110001"; z_correct<="0001101011011001";
        when 10546 => y_in <= "10101001"; x_in <= "10110010"; z_correct<="0001101010000010";
        when 10547 => y_in <= "10101001"; x_in <= "10110011"; z_correct<="0001101000101011";
        when 10548 => y_in <= "10101001"; x_in <= "10110100"; z_correct<="0001100111010100";
        when 10549 => y_in <= "10101001"; x_in <= "10110101"; z_correct<="0001100101111101";
        when 10550 => y_in <= "10101001"; x_in <= "10110110"; z_correct<="0001100100100110";
        when 10551 => y_in <= "10101001"; x_in <= "10110111"; z_correct<="0001100011001111";
        when 10552 => y_in <= "10101001"; x_in <= "10111000"; z_correct<="0001100001111000";
        when 10553 => y_in <= "10101001"; x_in <= "10111001"; z_correct<="0001100000100001";
        when 10554 => y_in <= "10101001"; x_in <= "10111010"; z_correct<="0001011111001010";
        when 10555 => y_in <= "10101001"; x_in <= "10111011"; z_correct<="0001011101110011";
        when 10556 => y_in <= "10101001"; x_in <= "10111100"; z_correct<="0001011100011100";
        when 10557 => y_in <= "10101001"; x_in <= "10111101"; z_correct<="0001011011000101";
        when 10558 => y_in <= "10101001"; x_in <= "10111110"; z_correct<="0001011001101110";
        when 10559 => y_in <= "10101001"; x_in <= "10111111"; z_correct<="0001011000010111";
        when 10560 => y_in <= "10101001"; x_in <= "11000000"; z_correct<="0001010111000000";
        when 10561 => y_in <= "10101001"; x_in <= "11000001"; z_correct<="0001010101101001";
        when 10562 => y_in <= "10101001"; x_in <= "11000010"; z_correct<="0001010100010010";
        when 10563 => y_in <= "10101001"; x_in <= "11000011"; z_correct<="0001010010111011";
        when 10564 => y_in <= "10101001"; x_in <= "11000100"; z_correct<="0001010001100100";
        when 10565 => y_in <= "10101001"; x_in <= "11000101"; z_correct<="0001010000001101";
        when 10566 => y_in <= "10101001"; x_in <= "11000110"; z_correct<="0001001110110110";
        when 10567 => y_in <= "10101001"; x_in <= "11000111"; z_correct<="0001001101011111";
        when 10568 => y_in <= "10101001"; x_in <= "11001000"; z_correct<="0001001100001000";
        when 10569 => y_in <= "10101001"; x_in <= "11001001"; z_correct<="0001001010110001";
        when 10570 => y_in <= "10101001"; x_in <= "11001010"; z_correct<="0001001001011010";
        when 10571 => y_in <= "10101001"; x_in <= "11001011"; z_correct<="0001001000000011";
        when 10572 => y_in <= "10101001"; x_in <= "11001100"; z_correct<="0001000110101100";
        when 10573 => y_in <= "10101001"; x_in <= "11001101"; z_correct<="0001000101010101";
        when 10574 => y_in <= "10101001"; x_in <= "11001110"; z_correct<="0001000011111110";
        when 10575 => y_in <= "10101001"; x_in <= "11001111"; z_correct<="0001000010100111";
        when 10576 => y_in <= "10101001"; x_in <= "11010000"; z_correct<="0001000001010000";
        when 10577 => y_in <= "10101001"; x_in <= "11010001"; z_correct<="0000111111111001";
        when 10578 => y_in <= "10101001"; x_in <= "11010010"; z_correct<="0000111110100010";
        when 10579 => y_in <= "10101001"; x_in <= "11010011"; z_correct<="0000111101001011";
        when 10580 => y_in <= "10101001"; x_in <= "11010100"; z_correct<="0000111011110100";
        when 10581 => y_in <= "10101001"; x_in <= "11010101"; z_correct<="0000111010011101";
        when 10582 => y_in <= "10101001"; x_in <= "11010110"; z_correct<="0000111001000110";
        when 10583 => y_in <= "10101001"; x_in <= "11010111"; z_correct<="0000110111101111";
        when 10584 => y_in <= "10101001"; x_in <= "11011000"; z_correct<="0000110110011000";
        when 10585 => y_in <= "10101001"; x_in <= "11011001"; z_correct<="0000110101000001";
        when 10586 => y_in <= "10101001"; x_in <= "11011010"; z_correct<="0000110011101010";
        when 10587 => y_in <= "10101001"; x_in <= "11011011"; z_correct<="0000110010010011";
        when 10588 => y_in <= "10101001"; x_in <= "11011100"; z_correct<="0000110000111100";
        when 10589 => y_in <= "10101001"; x_in <= "11011101"; z_correct<="0000101111100101";
        when 10590 => y_in <= "10101001"; x_in <= "11011110"; z_correct<="0000101110001110";
        when 10591 => y_in <= "10101001"; x_in <= "11011111"; z_correct<="0000101100110111";
        when 10592 => y_in <= "10101001"; x_in <= "11100000"; z_correct<="0000101011100000";
        when 10593 => y_in <= "10101001"; x_in <= "11100001"; z_correct<="0000101010001001";
        when 10594 => y_in <= "10101001"; x_in <= "11100010"; z_correct<="0000101000110010";
        when 10595 => y_in <= "10101001"; x_in <= "11100011"; z_correct<="0000100111011011";
        when 10596 => y_in <= "10101001"; x_in <= "11100100"; z_correct<="0000100110000100";
        when 10597 => y_in <= "10101001"; x_in <= "11100101"; z_correct<="0000100100101101";
        when 10598 => y_in <= "10101001"; x_in <= "11100110"; z_correct<="0000100011010110";
        when 10599 => y_in <= "10101001"; x_in <= "11100111"; z_correct<="0000100001111111";
        when 10600 => y_in <= "10101001"; x_in <= "11101000"; z_correct<="0000100000101000";
        when 10601 => y_in <= "10101001"; x_in <= "11101001"; z_correct<="0000011111010001";
        when 10602 => y_in <= "10101001"; x_in <= "11101010"; z_correct<="0000011101111010";
        when 10603 => y_in <= "10101001"; x_in <= "11101011"; z_correct<="0000011100100011";
        when 10604 => y_in <= "10101001"; x_in <= "11101100"; z_correct<="0000011011001100";
        when 10605 => y_in <= "10101001"; x_in <= "11101101"; z_correct<="0000011001110101";
        when 10606 => y_in <= "10101001"; x_in <= "11101110"; z_correct<="0000011000011110";
        when 10607 => y_in <= "10101001"; x_in <= "11101111"; z_correct<="0000010111000111";
        when 10608 => y_in <= "10101001"; x_in <= "11110000"; z_correct<="0000010101110000";
        when 10609 => y_in <= "10101001"; x_in <= "11110001"; z_correct<="0000010100011001";
        when 10610 => y_in <= "10101001"; x_in <= "11110010"; z_correct<="0000010011000010";
        when 10611 => y_in <= "10101001"; x_in <= "11110011"; z_correct<="0000010001101011";
        when 10612 => y_in <= "10101001"; x_in <= "11110100"; z_correct<="0000010000010100";
        when 10613 => y_in <= "10101001"; x_in <= "11110101"; z_correct<="0000001110111101";
        when 10614 => y_in <= "10101001"; x_in <= "11110110"; z_correct<="0000001101100110";
        when 10615 => y_in <= "10101001"; x_in <= "11110111"; z_correct<="0000001100001111";
        when 10616 => y_in <= "10101001"; x_in <= "11111000"; z_correct<="0000001010111000";
        when 10617 => y_in <= "10101001"; x_in <= "11111001"; z_correct<="0000001001100001";
        when 10618 => y_in <= "10101001"; x_in <= "11111010"; z_correct<="0000001000001010";
        when 10619 => y_in <= "10101001"; x_in <= "11111011"; z_correct<="0000000110110011";
        when 10620 => y_in <= "10101001"; x_in <= "11111100"; z_correct<="0000000101011100";
        when 10621 => y_in <= "10101001"; x_in <= "11111101"; z_correct<="0000000100000101";
        when 10622 => y_in <= "10101001"; x_in <= "11111110"; z_correct<="0000000010101110";
        when 10623 => y_in <= "10101001"; x_in <= "11111111"; z_correct<="0000000001010111";
        when 10624 => y_in <= "10101001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 10625 => y_in <= "10101001"; x_in <= "00000001"; z_correct<="1111111110101001";
        when 10626 => y_in <= "10101001"; x_in <= "00000010"; z_correct<="1111111101010010";
        when 10627 => y_in <= "10101001"; x_in <= "00000011"; z_correct<="1111111011111011";
        when 10628 => y_in <= "10101001"; x_in <= "00000100"; z_correct<="1111111010100100";
        when 10629 => y_in <= "10101001"; x_in <= "00000101"; z_correct<="1111111001001101";
        when 10630 => y_in <= "10101001"; x_in <= "00000110"; z_correct<="1111110111110110";
        when 10631 => y_in <= "10101001"; x_in <= "00000111"; z_correct<="1111110110011111";
        when 10632 => y_in <= "10101001"; x_in <= "00001000"; z_correct<="1111110101001000";
        when 10633 => y_in <= "10101001"; x_in <= "00001001"; z_correct<="1111110011110001";
        when 10634 => y_in <= "10101001"; x_in <= "00001010"; z_correct<="1111110010011010";
        when 10635 => y_in <= "10101001"; x_in <= "00001011"; z_correct<="1111110001000011";
        when 10636 => y_in <= "10101001"; x_in <= "00001100"; z_correct<="1111101111101100";
        when 10637 => y_in <= "10101001"; x_in <= "00001101"; z_correct<="1111101110010101";
        when 10638 => y_in <= "10101001"; x_in <= "00001110"; z_correct<="1111101100111110";
        when 10639 => y_in <= "10101001"; x_in <= "00001111"; z_correct<="1111101011100111";
        when 10640 => y_in <= "10101001"; x_in <= "00010000"; z_correct<="1111101010010000";
        when 10641 => y_in <= "10101001"; x_in <= "00010001"; z_correct<="1111101000111001";
        when 10642 => y_in <= "10101001"; x_in <= "00010010"; z_correct<="1111100111100010";
        when 10643 => y_in <= "10101001"; x_in <= "00010011"; z_correct<="1111100110001011";
        when 10644 => y_in <= "10101001"; x_in <= "00010100"; z_correct<="1111100100110100";
        when 10645 => y_in <= "10101001"; x_in <= "00010101"; z_correct<="1111100011011101";
        when 10646 => y_in <= "10101001"; x_in <= "00010110"; z_correct<="1111100010000110";
        when 10647 => y_in <= "10101001"; x_in <= "00010111"; z_correct<="1111100000101111";
        when 10648 => y_in <= "10101001"; x_in <= "00011000"; z_correct<="1111011111011000";
        when 10649 => y_in <= "10101001"; x_in <= "00011001"; z_correct<="1111011110000001";
        when 10650 => y_in <= "10101001"; x_in <= "00011010"; z_correct<="1111011100101010";
        when 10651 => y_in <= "10101001"; x_in <= "00011011"; z_correct<="1111011011010011";
        when 10652 => y_in <= "10101001"; x_in <= "00011100"; z_correct<="1111011001111100";
        when 10653 => y_in <= "10101001"; x_in <= "00011101"; z_correct<="1111011000100101";
        when 10654 => y_in <= "10101001"; x_in <= "00011110"; z_correct<="1111010111001110";
        when 10655 => y_in <= "10101001"; x_in <= "00011111"; z_correct<="1111010101110111";
        when 10656 => y_in <= "10101001"; x_in <= "00100000"; z_correct<="1111010100100000";
        when 10657 => y_in <= "10101001"; x_in <= "00100001"; z_correct<="1111010011001001";
        when 10658 => y_in <= "10101001"; x_in <= "00100010"; z_correct<="1111010001110010";
        when 10659 => y_in <= "10101001"; x_in <= "00100011"; z_correct<="1111010000011011";
        when 10660 => y_in <= "10101001"; x_in <= "00100100"; z_correct<="1111001111000100";
        when 10661 => y_in <= "10101001"; x_in <= "00100101"; z_correct<="1111001101101101";
        when 10662 => y_in <= "10101001"; x_in <= "00100110"; z_correct<="1111001100010110";
        when 10663 => y_in <= "10101001"; x_in <= "00100111"; z_correct<="1111001010111111";
        when 10664 => y_in <= "10101001"; x_in <= "00101000"; z_correct<="1111001001101000";
        when 10665 => y_in <= "10101001"; x_in <= "00101001"; z_correct<="1111001000010001";
        when 10666 => y_in <= "10101001"; x_in <= "00101010"; z_correct<="1111000110111010";
        when 10667 => y_in <= "10101001"; x_in <= "00101011"; z_correct<="1111000101100011";
        when 10668 => y_in <= "10101001"; x_in <= "00101100"; z_correct<="1111000100001100";
        when 10669 => y_in <= "10101001"; x_in <= "00101101"; z_correct<="1111000010110101";
        when 10670 => y_in <= "10101001"; x_in <= "00101110"; z_correct<="1111000001011110";
        when 10671 => y_in <= "10101001"; x_in <= "00101111"; z_correct<="1111000000000111";
        when 10672 => y_in <= "10101001"; x_in <= "00110000"; z_correct<="1110111110110000";
        when 10673 => y_in <= "10101001"; x_in <= "00110001"; z_correct<="1110111101011001";
        when 10674 => y_in <= "10101001"; x_in <= "00110010"; z_correct<="1110111100000010";
        when 10675 => y_in <= "10101001"; x_in <= "00110011"; z_correct<="1110111010101011";
        when 10676 => y_in <= "10101001"; x_in <= "00110100"; z_correct<="1110111001010100";
        when 10677 => y_in <= "10101001"; x_in <= "00110101"; z_correct<="1110110111111101";
        when 10678 => y_in <= "10101001"; x_in <= "00110110"; z_correct<="1110110110100110";
        when 10679 => y_in <= "10101001"; x_in <= "00110111"; z_correct<="1110110101001111";
        when 10680 => y_in <= "10101001"; x_in <= "00111000"; z_correct<="1110110011111000";
        when 10681 => y_in <= "10101001"; x_in <= "00111001"; z_correct<="1110110010100001";
        when 10682 => y_in <= "10101001"; x_in <= "00111010"; z_correct<="1110110001001010";
        when 10683 => y_in <= "10101001"; x_in <= "00111011"; z_correct<="1110101111110011";
        when 10684 => y_in <= "10101001"; x_in <= "00111100"; z_correct<="1110101110011100";
        when 10685 => y_in <= "10101001"; x_in <= "00111101"; z_correct<="1110101101000101";
        when 10686 => y_in <= "10101001"; x_in <= "00111110"; z_correct<="1110101011101110";
        when 10687 => y_in <= "10101001"; x_in <= "00111111"; z_correct<="1110101010010111";
        when 10688 => y_in <= "10101001"; x_in <= "01000000"; z_correct<="1110101001000000";
        when 10689 => y_in <= "10101001"; x_in <= "01000001"; z_correct<="1110100111101001";
        when 10690 => y_in <= "10101001"; x_in <= "01000010"; z_correct<="1110100110010010";
        when 10691 => y_in <= "10101001"; x_in <= "01000011"; z_correct<="1110100100111011";
        when 10692 => y_in <= "10101001"; x_in <= "01000100"; z_correct<="1110100011100100";
        when 10693 => y_in <= "10101001"; x_in <= "01000101"; z_correct<="1110100010001101";
        when 10694 => y_in <= "10101001"; x_in <= "01000110"; z_correct<="1110100000110110";
        when 10695 => y_in <= "10101001"; x_in <= "01000111"; z_correct<="1110011111011111";
        when 10696 => y_in <= "10101001"; x_in <= "01001000"; z_correct<="1110011110001000";
        when 10697 => y_in <= "10101001"; x_in <= "01001001"; z_correct<="1110011100110001";
        when 10698 => y_in <= "10101001"; x_in <= "01001010"; z_correct<="1110011011011010";
        when 10699 => y_in <= "10101001"; x_in <= "01001011"; z_correct<="1110011010000011";
        when 10700 => y_in <= "10101001"; x_in <= "01001100"; z_correct<="1110011000101100";
        when 10701 => y_in <= "10101001"; x_in <= "01001101"; z_correct<="1110010111010101";
        when 10702 => y_in <= "10101001"; x_in <= "01001110"; z_correct<="1110010101111110";
        when 10703 => y_in <= "10101001"; x_in <= "01001111"; z_correct<="1110010100100111";
        when 10704 => y_in <= "10101001"; x_in <= "01010000"; z_correct<="1110010011010000";
        when 10705 => y_in <= "10101001"; x_in <= "01010001"; z_correct<="1110010001111001";
        when 10706 => y_in <= "10101001"; x_in <= "01010010"; z_correct<="1110010000100010";
        when 10707 => y_in <= "10101001"; x_in <= "01010011"; z_correct<="1110001111001011";
        when 10708 => y_in <= "10101001"; x_in <= "01010100"; z_correct<="1110001101110100";
        when 10709 => y_in <= "10101001"; x_in <= "01010101"; z_correct<="1110001100011101";
        when 10710 => y_in <= "10101001"; x_in <= "01010110"; z_correct<="1110001011000110";
        when 10711 => y_in <= "10101001"; x_in <= "01010111"; z_correct<="1110001001101111";
        when 10712 => y_in <= "10101001"; x_in <= "01011000"; z_correct<="1110001000011000";
        when 10713 => y_in <= "10101001"; x_in <= "01011001"; z_correct<="1110000111000001";
        when 10714 => y_in <= "10101001"; x_in <= "01011010"; z_correct<="1110000101101010";
        when 10715 => y_in <= "10101001"; x_in <= "01011011"; z_correct<="1110000100010011";
        when 10716 => y_in <= "10101001"; x_in <= "01011100"; z_correct<="1110000010111100";
        when 10717 => y_in <= "10101001"; x_in <= "01011101"; z_correct<="1110000001100101";
        when 10718 => y_in <= "10101001"; x_in <= "01011110"; z_correct<="1110000000001110";
        when 10719 => y_in <= "10101001"; x_in <= "01011111"; z_correct<="1101111110110111";
        when 10720 => y_in <= "10101001"; x_in <= "01100000"; z_correct<="1101111101100000";
        when 10721 => y_in <= "10101001"; x_in <= "01100001"; z_correct<="1101111100001001";
        when 10722 => y_in <= "10101001"; x_in <= "01100010"; z_correct<="1101111010110010";
        when 10723 => y_in <= "10101001"; x_in <= "01100011"; z_correct<="1101111001011011";
        when 10724 => y_in <= "10101001"; x_in <= "01100100"; z_correct<="1101111000000100";
        when 10725 => y_in <= "10101001"; x_in <= "01100101"; z_correct<="1101110110101101";
        when 10726 => y_in <= "10101001"; x_in <= "01100110"; z_correct<="1101110101010110";
        when 10727 => y_in <= "10101001"; x_in <= "01100111"; z_correct<="1101110011111111";
        when 10728 => y_in <= "10101001"; x_in <= "01101000"; z_correct<="1101110010101000";
        when 10729 => y_in <= "10101001"; x_in <= "01101001"; z_correct<="1101110001010001";
        when 10730 => y_in <= "10101001"; x_in <= "01101010"; z_correct<="1101101111111010";
        when 10731 => y_in <= "10101001"; x_in <= "01101011"; z_correct<="1101101110100011";
        when 10732 => y_in <= "10101001"; x_in <= "01101100"; z_correct<="1101101101001100";
        when 10733 => y_in <= "10101001"; x_in <= "01101101"; z_correct<="1101101011110101";
        when 10734 => y_in <= "10101001"; x_in <= "01101110"; z_correct<="1101101010011110";
        when 10735 => y_in <= "10101001"; x_in <= "01101111"; z_correct<="1101101001000111";
        when 10736 => y_in <= "10101001"; x_in <= "01110000"; z_correct<="1101100111110000";
        when 10737 => y_in <= "10101001"; x_in <= "01110001"; z_correct<="1101100110011001";
        when 10738 => y_in <= "10101001"; x_in <= "01110010"; z_correct<="1101100101000010";
        when 10739 => y_in <= "10101001"; x_in <= "01110011"; z_correct<="1101100011101011";
        when 10740 => y_in <= "10101001"; x_in <= "01110100"; z_correct<="1101100010010100";
        when 10741 => y_in <= "10101001"; x_in <= "01110101"; z_correct<="1101100000111101";
        when 10742 => y_in <= "10101001"; x_in <= "01110110"; z_correct<="1101011111100110";
        when 10743 => y_in <= "10101001"; x_in <= "01110111"; z_correct<="1101011110001111";
        when 10744 => y_in <= "10101001"; x_in <= "01111000"; z_correct<="1101011100111000";
        when 10745 => y_in <= "10101001"; x_in <= "01111001"; z_correct<="1101011011100001";
        when 10746 => y_in <= "10101001"; x_in <= "01111010"; z_correct<="1101011010001010";
        when 10747 => y_in <= "10101001"; x_in <= "01111011"; z_correct<="1101011000110011";
        when 10748 => y_in <= "10101001"; x_in <= "01111100"; z_correct<="1101010111011100";
        when 10749 => y_in <= "10101001"; x_in <= "01111101"; z_correct<="1101010110000101";
        when 10750 => y_in <= "10101001"; x_in <= "01111110"; z_correct<="1101010100101110";
        when 10751 => y_in <= "10101001"; x_in <= "01111111"; z_correct<="1101010011010111";
        when 10752 => y_in <= "10101010"; x_in <= "10000000"; z_correct<="0010101100000000";
        when 10753 => y_in <= "10101010"; x_in <= "10000001"; z_correct<="0010101010101010";
        when 10754 => y_in <= "10101010"; x_in <= "10000010"; z_correct<="0010101001010100";
        when 10755 => y_in <= "10101010"; x_in <= "10000011"; z_correct<="0010100111111110";
        when 10756 => y_in <= "10101010"; x_in <= "10000100"; z_correct<="0010100110101000";
        when 10757 => y_in <= "10101010"; x_in <= "10000101"; z_correct<="0010100101010010";
        when 10758 => y_in <= "10101010"; x_in <= "10000110"; z_correct<="0010100011111100";
        when 10759 => y_in <= "10101010"; x_in <= "10000111"; z_correct<="0010100010100110";
        when 10760 => y_in <= "10101010"; x_in <= "10001000"; z_correct<="0010100001010000";
        when 10761 => y_in <= "10101010"; x_in <= "10001001"; z_correct<="0010011111111010";
        when 10762 => y_in <= "10101010"; x_in <= "10001010"; z_correct<="0010011110100100";
        when 10763 => y_in <= "10101010"; x_in <= "10001011"; z_correct<="0010011101001110";
        when 10764 => y_in <= "10101010"; x_in <= "10001100"; z_correct<="0010011011111000";
        when 10765 => y_in <= "10101010"; x_in <= "10001101"; z_correct<="0010011010100010";
        when 10766 => y_in <= "10101010"; x_in <= "10001110"; z_correct<="0010011001001100";
        when 10767 => y_in <= "10101010"; x_in <= "10001111"; z_correct<="0010010111110110";
        when 10768 => y_in <= "10101010"; x_in <= "10010000"; z_correct<="0010010110100000";
        when 10769 => y_in <= "10101010"; x_in <= "10010001"; z_correct<="0010010101001010";
        when 10770 => y_in <= "10101010"; x_in <= "10010010"; z_correct<="0010010011110100";
        when 10771 => y_in <= "10101010"; x_in <= "10010011"; z_correct<="0010010010011110";
        when 10772 => y_in <= "10101010"; x_in <= "10010100"; z_correct<="0010010001001000";
        when 10773 => y_in <= "10101010"; x_in <= "10010101"; z_correct<="0010001111110010";
        when 10774 => y_in <= "10101010"; x_in <= "10010110"; z_correct<="0010001110011100";
        when 10775 => y_in <= "10101010"; x_in <= "10010111"; z_correct<="0010001101000110";
        when 10776 => y_in <= "10101010"; x_in <= "10011000"; z_correct<="0010001011110000";
        when 10777 => y_in <= "10101010"; x_in <= "10011001"; z_correct<="0010001010011010";
        when 10778 => y_in <= "10101010"; x_in <= "10011010"; z_correct<="0010001001000100";
        when 10779 => y_in <= "10101010"; x_in <= "10011011"; z_correct<="0010000111101110";
        when 10780 => y_in <= "10101010"; x_in <= "10011100"; z_correct<="0010000110011000";
        when 10781 => y_in <= "10101010"; x_in <= "10011101"; z_correct<="0010000101000010";
        when 10782 => y_in <= "10101010"; x_in <= "10011110"; z_correct<="0010000011101100";
        when 10783 => y_in <= "10101010"; x_in <= "10011111"; z_correct<="0010000010010110";
        when 10784 => y_in <= "10101010"; x_in <= "10100000"; z_correct<="0010000001000000";
        when 10785 => y_in <= "10101010"; x_in <= "10100001"; z_correct<="0001111111101010";
        when 10786 => y_in <= "10101010"; x_in <= "10100010"; z_correct<="0001111110010100";
        when 10787 => y_in <= "10101010"; x_in <= "10100011"; z_correct<="0001111100111110";
        when 10788 => y_in <= "10101010"; x_in <= "10100100"; z_correct<="0001111011101000";
        when 10789 => y_in <= "10101010"; x_in <= "10100101"; z_correct<="0001111010010010";
        when 10790 => y_in <= "10101010"; x_in <= "10100110"; z_correct<="0001111000111100";
        when 10791 => y_in <= "10101010"; x_in <= "10100111"; z_correct<="0001110111100110";
        when 10792 => y_in <= "10101010"; x_in <= "10101000"; z_correct<="0001110110010000";
        when 10793 => y_in <= "10101010"; x_in <= "10101001"; z_correct<="0001110100111010";
        when 10794 => y_in <= "10101010"; x_in <= "10101010"; z_correct<="0001110011100100";
        when 10795 => y_in <= "10101010"; x_in <= "10101011"; z_correct<="0001110010001110";
        when 10796 => y_in <= "10101010"; x_in <= "10101100"; z_correct<="0001110000111000";
        when 10797 => y_in <= "10101010"; x_in <= "10101101"; z_correct<="0001101111100010";
        when 10798 => y_in <= "10101010"; x_in <= "10101110"; z_correct<="0001101110001100";
        when 10799 => y_in <= "10101010"; x_in <= "10101111"; z_correct<="0001101100110110";
        when 10800 => y_in <= "10101010"; x_in <= "10110000"; z_correct<="0001101011100000";
        when 10801 => y_in <= "10101010"; x_in <= "10110001"; z_correct<="0001101010001010";
        when 10802 => y_in <= "10101010"; x_in <= "10110010"; z_correct<="0001101000110100";
        when 10803 => y_in <= "10101010"; x_in <= "10110011"; z_correct<="0001100111011110";
        when 10804 => y_in <= "10101010"; x_in <= "10110100"; z_correct<="0001100110001000";
        when 10805 => y_in <= "10101010"; x_in <= "10110101"; z_correct<="0001100100110010";
        when 10806 => y_in <= "10101010"; x_in <= "10110110"; z_correct<="0001100011011100";
        when 10807 => y_in <= "10101010"; x_in <= "10110111"; z_correct<="0001100010000110";
        when 10808 => y_in <= "10101010"; x_in <= "10111000"; z_correct<="0001100000110000";
        when 10809 => y_in <= "10101010"; x_in <= "10111001"; z_correct<="0001011111011010";
        when 10810 => y_in <= "10101010"; x_in <= "10111010"; z_correct<="0001011110000100";
        when 10811 => y_in <= "10101010"; x_in <= "10111011"; z_correct<="0001011100101110";
        when 10812 => y_in <= "10101010"; x_in <= "10111100"; z_correct<="0001011011011000";
        when 10813 => y_in <= "10101010"; x_in <= "10111101"; z_correct<="0001011010000010";
        when 10814 => y_in <= "10101010"; x_in <= "10111110"; z_correct<="0001011000101100";
        when 10815 => y_in <= "10101010"; x_in <= "10111111"; z_correct<="0001010111010110";
        when 10816 => y_in <= "10101010"; x_in <= "11000000"; z_correct<="0001010110000000";
        when 10817 => y_in <= "10101010"; x_in <= "11000001"; z_correct<="0001010100101010";
        when 10818 => y_in <= "10101010"; x_in <= "11000010"; z_correct<="0001010011010100";
        when 10819 => y_in <= "10101010"; x_in <= "11000011"; z_correct<="0001010001111110";
        when 10820 => y_in <= "10101010"; x_in <= "11000100"; z_correct<="0001010000101000";
        when 10821 => y_in <= "10101010"; x_in <= "11000101"; z_correct<="0001001111010010";
        when 10822 => y_in <= "10101010"; x_in <= "11000110"; z_correct<="0001001101111100";
        when 10823 => y_in <= "10101010"; x_in <= "11000111"; z_correct<="0001001100100110";
        when 10824 => y_in <= "10101010"; x_in <= "11001000"; z_correct<="0001001011010000";
        when 10825 => y_in <= "10101010"; x_in <= "11001001"; z_correct<="0001001001111010";
        when 10826 => y_in <= "10101010"; x_in <= "11001010"; z_correct<="0001001000100100";
        when 10827 => y_in <= "10101010"; x_in <= "11001011"; z_correct<="0001000111001110";
        when 10828 => y_in <= "10101010"; x_in <= "11001100"; z_correct<="0001000101111000";
        when 10829 => y_in <= "10101010"; x_in <= "11001101"; z_correct<="0001000100100010";
        when 10830 => y_in <= "10101010"; x_in <= "11001110"; z_correct<="0001000011001100";
        when 10831 => y_in <= "10101010"; x_in <= "11001111"; z_correct<="0001000001110110";
        when 10832 => y_in <= "10101010"; x_in <= "11010000"; z_correct<="0001000000100000";
        when 10833 => y_in <= "10101010"; x_in <= "11010001"; z_correct<="0000111111001010";
        when 10834 => y_in <= "10101010"; x_in <= "11010010"; z_correct<="0000111101110100";
        when 10835 => y_in <= "10101010"; x_in <= "11010011"; z_correct<="0000111100011110";
        when 10836 => y_in <= "10101010"; x_in <= "11010100"; z_correct<="0000111011001000";
        when 10837 => y_in <= "10101010"; x_in <= "11010101"; z_correct<="0000111001110010";
        when 10838 => y_in <= "10101010"; x_in <= "11010110"; z_correct<="0000111000011100";
        when 10839 => y_in <= "10101010"; x_in <= "11010111"; z_correct<="0000110111000110";
        when 10840 => y_in <= "10101010"; x_in <= "11011000"; z_correct<="0000110101110000";
        when 10841 => y_in <= "10101010"; x_in <= "11011001"; z_correct<="0000110100011010";
        when 10842 => y_in <= "10101010"; x_in <= "11011010"; z_correct<="0000110011000100";
        when 10843 => y_in <= "10101010"; x_in <= "11011011"; z_correct<="0000110001101110";
        when 10844 => y_in <= "10101010"; x_in <= "11011100"; z_correct<="0000110000011000";
        when 10845 => y_in <= "10101010"; x_in <= "11011101"; z_correct<="0000101111000010";
        when 10846 => y_in <= "10101010"; x_in <= "11011110"; z_correct<="0000101101101100";
        when 10847 => y_in <= "10101010"; x_in <= "11011111"; z_correct<="0000101100010110";
        when 10848 => y_in <= "10101010"; x_in <= "11100000"; z_correct<="0000101011000000";
        when 10849 => y_in <= "10101010"; x_in <= "11100001"; z_correct<="0000101001101010";
        when 10850 => y_in <= "10101010"; x_in <= "11100010"; z_correct<="0000101000010100";
        when 10851 => y_in <= "10101010"; x_in <= "11100011"; z_correct<="0000100110111110";
        when 10852 => y_in <= "10101010"; x_in <= "11100100"; z_correct<="0000100101101000";
        when 10853 => y_in <= "10101010"; x_in <= "11100101"; z_correct<="0000100100010010";
        when 10854 => y_in <= "10101010"; x_in <= "11100110"; z_correct<="0000100010111100";
        when 10855 => y_in <= "10101010"; x_in <= "11100111"; z_correct<="0000100001100110";
        when 10856 => y_in <= "10101010"; x_in <= "11101000"; z_correct<="0000100000010000";
        when 10857 => y_in <= "10101010"; x_in <= "11101001"; z_correct<="0000011110111010";
        when 10858 => y_in <= "10101010"; x_in <= "11101010"; z_correct<="0000011101100100";
        when 10859 => y_in <= "10101010"; x_in <= "11101011"; z_correct<="0000011100001110";
        when 10860 => y_in <= "10101010"; x_in <= "11101100"; z_correct<="0000011010111000";
        when 10861 => y_in <= "10101010"; x_in <= "11101101"; z_correct<="0000011001100010";
        when 10862 => y_in <= "10101010"; x_in <= "11101110"; z_correct<="0000011000001100";
        when 10863 => y_in <= "10101010"; x_in <= "11101111"; z_correct<="0000010110110110";
        when 10864 => y_in <= "10101010"; x_in <= "11110000"; z_correct<="0000010101100000";
        when 10865 => y_in <= "10101010"; x_in <= "11110001"; z_correct<="0000010100001010";
        when 10866 => y_in <= "10101010"; x_in <= "11110010"; z_correct<="0000010010110100";
        when 10867 => y_in <= "10101010"; x_in <= "11110011"; z_correct<="0000010001011110";
        when 10868 => y_in <= "10101010"; x_in <= "11110100"; z_correct<="0000010000001000";
        when 10869 => y_in <= "10101010"; x_in <= "11110101"; z_correct<="0000001110110010";
        when 10870 => y_in <= "10101010"; x_in <= "11110110"; z_correct<="0000001101011100";
        when 10871 => y_in <= "10101010"; x_in <= "11110111"; z_correct<="0000001100000110";
        when 10872 => y_in <= "10101010"; x_in <= "11111000"; z_correct<="0000001010110000";
        when 10873 => y_in <= "10101010"; x_in <= "11111001"; z_correct<="0000001001011010";
        when 10874 => y_in <= "10101010"; x_in <= "11111010"; z_correct<="0000001000000100";
        when 10875 => y_in <= "10101010"; x_in <= "11111011"; z_correct<="0000000110101110";
        when 10876 => y_in <= "10101010"; x_in <= "11111100"; z_correct<="0000000101011000";
        when 10877 => y_in <= "10101010"; x_in <= "11111101"; z_correct<="0000000100000010";
        when 10878 => y_in <= "10101010"; x_in <= "11111110"; z_correct<="0000000010101100";
        when 10879 => y_in <= "10101010"; x_in <= "11111111"; z_correct<="0000000001010110";
        when 10880 => y_in <= "10101010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 10881 => y_in <= "10101010"; x_in <= "00000001"; z_correct<="1111111110101010";
        when 10882 => y_in <= "10101010"; x_in <= "00000010"; z_correct<="1111111101010100";
        when 10883 => y_in <= "10101010"; x_in <= "00000011"; z_correct<="1111111011111110";
        when 10884 => y_in <= "10101010"; x_in <= "00000100"; z_correct<="1111111010101000";
        when 10885 => y_in <= "10101010"; x_in <= "00000101"; z_correct<="1111111001010010";
        when 10886 => y_in <= "10101010"; x_in <= "00000110"; z_correct<="1111110111111100";
        when 10887 => y_in <= "10101010"; x_in <= "00000111"; z_correct<="1111110110100110";
        when 10888 => y_in <= "10101010"; x_in <= "00001000"; z_correct<="1111110101010000";
        when 10889 => y_in <= "10101010"; x_in <= "00001001"; z_correct<="1111110011111010";
        when 10890 => y_in <= "10101010"; x_in <= "00001010"; z_correct<="1111110010100100";
        when 10891 => y_in <= "10101010"; x_in <= "00001011"; z_correct<="1111110001001110";
        when 10892 => y_in <= "10101010"; x_in <= "00001100"; z_correct<="1111101111111000";
        when 10893 => y_in <= "10101010"; x_in <= "00001101"; z_correct<="1111101110100010";
        when 10894 => y_in <= "10101010"; x_in <= "00001110"; z_correct<="1111101101001100";
        when 10895 => y_in <= "10101010"; x_in <= "00001111"; z_correct<="1111101011110110";
        when 10896 => y_in <= "10101010"; x_in <= "00010000"; z_correct<="1111101010100000";
        when 10897 => y_in <= "10101010"; x_in <= "00010001"; z_correct<="1111101001001010";
        when 10898 => y_in <= "10101010"; x_in <= "00010010"; z_correct<="1111100111110100";
        when 10899 => y_in <= "10101010"; x_in <= "00010011"; z_correct<="1111100110011110";
        when 10900 => y_in <= "10101010"; x_in <= "00010100"; z_correct<="1111100101001000";
        when 10901 => y_in <= "10101010"; x_in <= "00010101"; z_correct<="1111100011110010";
        when 10902 => y_in <= "10101010"; x_in <= "00010110"; z_correct<="1111100010011100";
        when 10903 => y_in <= "10101010"; x_in <= "00010111"; z_correct<="1111100001000110";
        when 10904 => y_in <= "10101010"; x_in <= "00011000"; z_correct<="1111011111110000";
        when 10905 => y_in <= "10101010"; x_in <= "00011001"; z_correct<="1111011110011010";
        when 10906 => y_in <= "10101010"; x_in <= "00011010"; z_correct<="1111011101000100";
        when 10907 => y_in <= "10101010"; x_in <= "00011011"; z_correct<="1111011011101110";
        when 10908 => y_in <= "10101010"; x_in <= "00011100"; z_correct<="1111011010011000";
        when 10909 => y_in <= "10101010"; x_in <= "00011101"; z_correct<="1111011001000010";
        when 10910 => y_in <= "10101010"; x_in <= "00011110"; z_correct<="1111010111101100";
        when 10911 => y_in <= "10101010"; x_in <= "00011111"; z_correct<="1111010110010110";
        when 10912 => y_in <= "10101010"; x_in <= "00100000"; z_correct<="1111010101000000";
        when 10913 => y_in <= "10101010"; x_in <= "00100001"; z_correct<="1111010011101010";
        when 10914 => y_in <= "10101010"; x_in <= "00100010"; z_correct<="1111010010010100";
        when 10915 => y_in <= "10101010"; x_in <= "00100011"; z_correct<="1111010000111110";
        when 10916 => y_in <= "10101010"; x_in <= "00100100"; z_correct<="1111001111101000";
        when 10917 => y_in <= "10101010"; x_in <= "00100101"; z_correct<="1111001110010010";
        when 10918 => y_in <= "10101010"; x_in <= "00100110"; z_correct<="1111001100111100";
        when 10919 => y_in <= "10101010"; x_in <= "00100111"; z_correct<="1111001011100110";
        when 10920 => y_in <= "10101010"; x_in <= "00101000"; z_correct<="1111001010010000";
        when 10921 => y_in <= "10101010"; x_in <= "00101001"; z_correct<="1111001000111010";
        when 10922 => y_in <= "10101010"; x_in <= "00101010"; z_correct<="1111000111100100";
        when 10923 => y_in <= "10101010"; x_in <= "00101011"; z_correct<="1111000110001110";
        when 10924 => y_in <= "10101010"; x_in <= "00101100"; z_correct<="1111000100111000";
        when 10925 => y_in <= "10101010"; x_in <= "00101101"; z_correct<="1111000011100010";
        when 10926 => y_in <= "10101010"; x_in <= "00101110"; z_correct<="1111000010001100";
        when 10927 => y_in <= "10101010"; x_in <= "00101111"; z_correct<="1111000000110110";
        when 10928 => y_in <= "10101010"; x_in <= "00110000"; z_correct<="1110111111100000";
        when 10929 => y_in <= "10101010"; x_in <= "00110001"; z_correct<="1110111110001010";
        when 10930 => y_in <= "10101010"; x_in <= "00110010"; z_correct<="1110111100110100";
        when 10931 => y_in <= "10101010"; x_in <= "00110011"; z_correct<="1110111011011110";
        when 10932 => y_in <= "10101010"; x_in <= "00110100"; z_correct<="1110111010001000";
        when 10933 => y_in <= "10101010"; x_in <= "00110101"; z_correct<="1110111000110010";
        when 10934 => y_in <= "10101010"; x_in <= "00110110"; z_correct<="1110110111011100";
        when 10935 => y_in <= "10101010"; x_in <= "00110111"; z_correct<="1110110110000110";
        when 10936 => y_in <= "10101010"; x_in <= "00111000"; z_correct<="1110110100110000";
        when 10937 => y_in <= "10101010"; x_in <= "00111001"; z_correct<="1110110011011010";
        when 10938 => y_in <= "10101010"; x_in <= "00111010"; z_correct<="1110110010000100";
        when 10939 => y_in <= "10101010"; x_in <= "00111011"; z_correct<="1110110000101110";
        when 10940 => y_in <= "10101010"; x_in <= "00111100"; z_correct<="1110101111011000";
        when 10941 => y_in <= "10101010"; x_in <= "00111101"; z_correct<="1110101110000010";
        when 10942 => y_in <= "10101010"; x_in <= "00111110"; z_correct<="1110101100101100";
        when 10943 => y_in <= "10101010"; x_in <= "00111111"; z_correct<="1110101011010110";
        when 10944 => y_in <= "10101010"; x_in <= "01000000"; z_correct<="1110101010000000";
        when 10945 => y_in <= "10101010"; x_in <= "01000001"; z_correct<="1110101000101010";
        when 10946 => y_in <= "10101010"; x_in <= "01000010"; z_correct<="1110100111010100";
        when 10947 => y_in <= "10101010"; x_in <= "01000011"; z_correct<="1110100101111110";
        when 10948 => y_in <= "10101010"; x_in <= "01000100"; z_correct<="1110100100101000";
        when 10949 => y_in <= "10101010"; x_in <= "01000101"; z_correct<="1110100011010010";
        when 10950 => y_in <= "10101010"; x_in <= "01000110"; z_correct<="1110100001111100";
        when 10951 => y_in <= "10101010"; x_in <= "01000111"; z_correct<="1110100000100110";
        when 10952 => y_in <= "10101010"; x_in <= "01001000"; z_correct<="1110011111010000";
        when 10953 => y_in <= "10101010"; x_in <= "01001001"; z_correct<="1110011101111010";
        when 10954 => y_in <= "10101010"; x_in <= "01001010"; z_correct<="1110011100100100";
        when 10955 => y_in <= "10101010"; x_in <= "01001011"; z_correct<="1110011011001110";
        when 10956 => y_in <= "10101010"; x_in <= "01001100"; z_correct<="1110011001111000";
        when 10957 => y_in <= "10101010"; x_in <= "01001101"; z_correct<="1110011000100010";
        when 10958 => y_in <= "10101010"; x_in <= "01001110"; z_correct<="1110010111001100";
        when 10959 => y_in <= "10101010"; x_in <= "01001111"; z_correct<="1110010101110110";
        when 10960 => y_in <= "10101010"; x_in <= "01010000"; z_correct<="1110010100100000";
        when 10961 => y_in <= "10101010"; x_in <= "01010001"; z_correct<="1110010011001010";
        when 10962 => y_in <= "10101010"; x_in <= "01010010"; z_correct<="1110010001110100";
        when 10963 => y_in <= "10101010"; x_in <= "01010011"; z_correct<="1110010000011110";
        when 10964 => y_in <= "10101010"; x_in <= "01010100"; z_correct<="1110001111001000";
        when 10965 => y_in <= "10101010"; x_in <= "01010101"; z_correct<="1110001101110010";
        when 10966 => y_in <= "10101010"; x_in <= "01010110"; z_correct<="1110001100011100";
        when 10967 => y_in <= "10101010"; x_in <= "01010111"; z_correct<="1110001011000110";
        when 10968 => y_in <= "10101010"; x_in <= "01011000"; z_correct<="1110001001110000";
        when 10969 => y_in <= "10101010"; x_in <= "01011001"; z_correct<="1110001000011010";
        when 10970 => y_in <= "10101010"; x_in <= "01011010"; z_correct<="1110000111000100";
        when 10971 => y_in <= "10101010"; x_in <= "01011011"; z_correct<="1110000101101110";
        when 10972 => y_in <= "10101010"; x_in <= "01011100"; z_correct<="1110000100011000";
        when 10973 => y_in <= "10101010"; x_in <= "01011101"; z_correct<="1110000011000010";
        when 10974 => y_in <= "10101010"; x_in <= "01011110"; z_correct<="1110000001101100";
        when 10975 => y_in <= "10101010"; x_in <= "01011111"; z_correct<="1110000000010110";
        when 10976 => y_in <= "10101010"; x_in <= "01100000"; z_correct<="1101111111000000";
        when 10977 => y_in <= "10101010"; x_in <= "01100001"; z_correct<="1101111101101010";
        when 10978 => y_in <= "10101010"; x_in <= "01100010"; z_correct<="1101111100010100";
        when 10979 => y_in <= "10101010"; x_in <= "01100011"; z_correct<="1101111010111110";
        when 10980 => y_in <= "10101010"; x_in <= "01100100"; z_correct<="1101111001101000";
        when 10981 => y_in <= "10101010"; x_in <= "01100101"; z_correct<="1101111000010010";
        when 10982 => y_in <= "10101010"; x_in <= "01100110"; z_correct<="1101110110111100";
        when 10983 => y_in <= "10101010"; x_in <= "01100111"; z_correct<="1101110101100110";
        when 10984 => y_in <= "10101010"; x_in <= "01101000"; z_correct<="1101110100010000";
        when 10985 => y_in <= "10101010"; x_in <= "01101001"; z_correct<="1101110010111010";
        when 10986 => y_in <= "10101010"; x_in <= "01101010"; z_correct<="1101110001100100";
        when 10987 => y_in <= "10101010"; x_in <= "01101011"; z_correct<="1101110000001110";
        when 10988 => y_in <= "10101010"; x_in <= "01101100"; z_correct<="1101101110111000";
        when 10989 => y_in <= "10101010"; x_in <= "01101101"; z_correct<="1101101101100010";
        when 10990 => y_in <= "10101010"; x_in <= "01101110"; z_correct<="1101101100001100";
        when 10991 => y_in <= "10101010"; x_in <= "01101111"; z_correct<="1101101010110110";
        when 10992 => y_in <= "10101010"; x_in <= "01110000"; z_correct<="1101101001100000";
        when 10993 => y_in <= "10101010"; x_in <= "01110001"; z_correct<="1101101000001010";
        when 10994 => y_in <= "10101010"; x_in <= "01110010"; z_correct<="1101100110110100";
        when 10995 => y_in <= "10101010"; x_in <= "01110011"; z_correct<="1101100101011110";
        when 10996 => y_in <= "10101010"; x_in <= "01110100"; z_correct<="1101100100001000";
        when 10997 => y_in <= "10101010"; x_in <= "01110101"; z_correct<="1101100010110010";
        when 10998 => y_in <= "10101010"; x_in <= "01110110"; z_correct<="1101100001011100";
        when 10999 => y_in <= "10101010"; x_in <= "01110111"; z_correct<="1101100000000110";
        when 11000 => y_in <= "10101010"; x_in <= "01111000"; z_correct<="1101011110110000";
        when 11001 => y_in <= "10101010"; x_in <= "01111001"; z_correct<="1101011101011010";
        when 11002 => y_in <= "10101010"; x_in <= "01111010"; z_correct<="1101011100000100";
        when 11003 => y_in <= "10101010"; x_in <= "01111011"; z_correct<="1101011010101110";
        when 11004 => y_in <= "10101010"; x_in <= "01111100"; z_correct<="1101011001011000";
        when 11005 => y_in <= "10101010"; x_in <= "01111101"; z_correct<="1101011000000010";
        when 11006 => y_in <= "10101010"; x_in <= "01111110"; z_correct<="1101010110101100";
        when 11007 => y_in <= "10101010"; x_in <= "01111111"; z_correct<="1101010101010110";
        when 11008 => y_in <= "10101011"; x_in <= "10000000"; z_correct<="0010101010000000";
        when 11009 => y_in <= "10101011"; x_in <= "10000001"; z_correct<="0010101000101011";
        when 11010 => y_in <= "10101011"; x_in <= "10000010"; z_correct<="0010100111010110";
        when 11011 => y_in <= "10101011"; x_in <= "10000011"; z_correct<="0010100110000001";
        when 11012 => y_in <= "10101011"; x_in <= "10000100"; z_correct<="0010100100101100";
        when 11013 => y_in <= "10101011"; x_in <= "10000101"; z_correct<="0010100011010111";
        when 11014 => y_in <= "10101011"; x_in <= "10000110"; z_correct<="0010100010000010";
        when 11015 => y_in <= "10101011"; x_in <= "10000111"; z_correct<="0010100000101101";
        when 11016 => y_in <= "10101011"; x_in <= "10001000"; z_correct<="0010011111011000";
        when 11017 => y_in <= "10101011"; x_in <= "10001001"; z_correct<="0010011110000011";
        when 11018 => y_in <= "10101011"; x_in <= "10001010"; z_correct<="0010011100101110";
        when 11019 => y_in <= "10101011"; x_in <= "10001011"; z_correct<="0010011011011001";
        when 11020 => y_in <= "10101011"; x_in <= "10001100"; z_correct<="0010011010000100";
        when 11021 => y_in <= "10101011"; x_in <= "10001101"; z_correct<="0010011000101111";
        when 11022 => y_in <= "10101011"; x_in <= "10001110"; z_correct<="0010010111011010";
        when 11023 => y_in <= "10101011"; x_in <= "10001111"; z_correct<="0010010110000101";
        when 11024 => y_in <= "10101011"; x_in <= "10010000"; z_correct<="0010010100110000";
        when 11025 => y_in <= "10101011"; x_in <= "10010001"; z_correct<="0010010011011011";
        when 11026 => y_in <= "10101011"; x_in <= "10010010"; z_correct<="0010010010000110";
        when 11027 => y_in <= "10101011"; x_in <= "10010011"; z_correct<="0010010000110001";
        when 11028 => y_in <= "10101011"; x_in <= "10010100"; z_correct<="0010001111011100";
        when 11029 => y_in <= "10101011"; x_in <= "10010101"; z_correct<="0010001110000111";
        when 11030 => y_in <= "10101011"; x_in <= "10010110"; z_correct<="0010001100110010";
        when 11031 => y_in <= "10101011"; x_in <= "10010111"; z_correct<="0010001011011101";
        when 11032 => y_in <= "10101011"; x_in <= "10011000"; z_correct<="0010001010001000";
        when 11033 => y_in <= "10101011"; x_in <= "10011001"; z_correct<="0010001000110011";
        when 11034 => y_in <= "10101011"; x_in <= "10011010"; z_correct<="0010000111011110";
        when 11035 => y_in <= "10101011"; x_in <= "10011011"; z_correct<="0010000110001001";
        when 11036 => y_in <= "10101011"; x_in <= "10011100"; z_correct<="0010000100110100";
        when 11037 => y_in <= "10101011"; x_in <= "10011101"; z_correct<="0010000011011111";
        when 11038 => y_in <= "10101011"; x_in <= "10011110"; z_correct<="0010000010001010";
        when 11039 => y_in <= "10101011"; x_in <= "10011111"; z_correct<="0010000000110101";
        when 11040 => y_in <= "10101011"; x_in <= "10100000"; z_correct<="0001111111100000";
        when 11041 => y_in <= "10101011"; x_in <= "10100001"; z_correct<="0001111110001011";
        when 11042 => y_in <= "10101011"; x_in <= "10100010"; z_correct<="0001111100110110";
        when 11043 => y_in <= "10101011"; x_in <= "10100011"; z_correct<="0001111011100001";
        when 11044 => y_in <= "10101011"; x_in <= "10100100"; z_correct<="0001111010001100";
        when 11045 => y_in <= "10101011"; x_in <= "10100101"; z_correct<="0001111000110111";
        when 11046 => y_in <= "10101011"; x_in <= "10100110"; z_correct<="0001110111100010";
        when 11047 => y_in <= "10101011"; x_in <= "10100111"; z_correct<="0001110110001101";
        when 11048 => y_in <= "10101011"; x_in <= "10101000"; z_correct<="0001110100111000";
        when 11049 => y_in <= "10101011"; x_in <= "10101001"; z_correct<="0001110011100011";
        when 11050 => y_in <= "10101011"; x_in <= "10101010"; z_correct<="0001110010001110";
        when 11051 => y_in <= "10101011"; x_in <= "10101011"; z_correct<="0001110000111001";
        when 11052 => y_in <= "10101011"; x_in <= "10101100"; z_correct<="0001101111100100";
        when 11053 => y_in <= "10101011"; x_in <= "10101101"; z_correct<="0001101110001111";
        when 11054 => y_in <= "10101011"; x_in <= "10101110"; z_correct<="0001101100111010";
        when 11055 => y_in <= "10101011"; x_in <= "10101111"; z_correct<="0001101011100101";
        when 11056 => y_in <= "10101011"; x_in <= "10110000"; z_correct<="0001101010010000";
        when 11057 => y_in <= "10101011"; x_in <= "10110001"; z_correct<="0001101000111011";
        when 11058 => y_in <= "10101011"; x_in <= "10110010"; z_correct<="0001100111100110";
        when 11059 => y_in <= "10101011"; x_in <= "10110011"; z_correct<="0001100110010001";
        when 11060 => y_in <= "10101011"; x_in <= "10110100"; z_correct<="0001100100111100";
        when 11061 => y_in <= "10101011"; x_in <= "10110101"; z_correct<="0001100011100111";
        when 11062 => y_in <= "10101011"; x_in <= "10110110"; z_correct<="0001100010010010";
        when 11063 => y_in <= "10101011"; x_in <= "10110111"; z_correct<="0001100000111101";
        when 11064 => y_in <= "10101011"; x_in <= "10111000"; z_correct<="0001011111101000";
        when 11065 => y_in <= "10101011"; x_in <= "10111001"; z_correct<="0001011110010011";
        when 11066 => y_in <= "10101011"; x_in <= "10111010"; z_correct<="0001011100111110";
        when 11067 => y_in <= "10101011"; x_in <= "10111011"; z_correct<="0001011011101001";
        when 11068 => y_in <= "10101011"; x_in <= "10111100"; z_correct<="0001011010010100";
        when 11069 => y_in <= "10101011"; x_in <= "10111101"; z_correct<="0001011000111111";
        when 11070 => y_in <= "10101011"; x_in <= "10111110"; z_correct<="0001010111101010";
        when 11071 => y_in <= "10101011"; x_in <= "10111111"; z_correct<="0001010110010101";
        when 11072 => y_in <= "10101011"; x_in <= "11000000"; z_correct<="0001010101000000";
        when 11073 => y_in <= "10101011"; x_in <= "11000001"; z_correct<="0001010011101011";
        when 11074 => y_in <= "10101011"; x_in <= "11000010"; z_correct<="0001010010010110";
        when 11075 => y_in <= "10101011"; x_in <= "11000011"; z_correct<="0001010001000001";
        when 11076 => y_in <= "10101011"; x_in <= "11000100"; z_correct<="0001001111101100";
        when 11077 => y_in <= "10101011"; x_in <= "11000101"; z_correct<="0001001110010111";
        when 11078 => y_in <= "10101011"; x_in <= "11000110"; z_correct<="0001001101000010";
        when 11079 => y_in <= "10101011"; x_in <= "11000111"; z_correct<="0001001011101101";
        when 11080 => y_in <= "10101011"; x_in <= "11001000"; z_correct<="0001001010011000";
        when 11081 => y_in <= "10101011"; x_in <= "11001001"; z_correct<="0001001001000011";
        when 11082 => y_in <= "10101011"; x_in <= "11001010"; z_correct<="0001000111101110";
        when 11083 => y_in <= "10101011"; x_in <= "11001011"; z_correct<="0001000110011001";
        when 11084 => y_in <= "10101011"; x_in <= "11001100"; z_correct<="0001000101000100";
        when 11085 => y_in <= "10101011"; x_in <= "11001101"; z_correct<="0001000011101111";
        when 11086 => y_in <= "10101011"; x_in <= "11001110"; z_correct<="0001000010011010";
        when 11087 => y_in <= "10101011"; x_in <= "11001111"; z_correct<="0001000001000101";
        when 11088 => y_in <= "10101011"; x_in <= "11010000"; z_correct<="0000111111110000";
        when 11089 => y_in <= "10101011"; x_in <= "11010001"; z_correct<="0000111110011011";
        when 11090 => y_in <= "10101011"; x_in <= "11010010"; z_correct<="0000111101000110";
        when 11091 => y_in <= "10101011"; x_in <= "11010011"; z_correct<="0000111011110001";
        when 11092 => y_in <= "10101011"; x_in <= "11010100"; z_correct<="0000111010011100";
        when 11093 => y_in <= "10101011"; x_in <= "11010101"; z_correct<="0000111001000111";
        when 11094 => y_in <= "10101011"; x_in <= "11010110"; z_correct<="0000110111110010";
        when 11095 => y_in <= "10101011"; x_in <= "11010111"; z_correct<="0000110110011101";
        when 11096 => y_in <= "10101011"; x_in <= "11011000"; z_correct<="0000110101001000";
        when 11097 => y_in <= "10101011"; x_in <= "11011001"; z_correct<="0000110011110011";
        when 11098 => y_in <= "10101011"; x_in <= "11011010"; z_correct<="0000110010011110";
        when 11099 => y_in <= "10101011"; x_in <= "11011011"; z_correct<="0000110001001001";
        when 11100 => y_in <= "10101011"; x_in <= "11011100"; z_correct<="0000101111110100";
        when 11101 => y_in <= "10101011"; x_in <= "11011101"; z_correct<="0000101110011111";
        when 11102 => y_in <= "10101011"; x_in <= "11011110"; z_correct<="0000101101001010";
        when 11103 => y_in <= "10101011"; x_in <= "11011111"; z_correct<="0000101011110101";
        when 11104 => y_in <= "10101011"; x_in <= "11100000"; z_correct<="0000101010100000";
        when 11105 => y_in <= "10101011"; x_in <= "11100001"; z_correct<="0000101001001011";
        when 11106 => y_in <= "10101011"; x_in <= "11100010"; z_correct<="0000100111110110";
        when 11107 => y_in <= "10101011"; x_in <= "11100011"; z_correct<="0000100110100001";
        when 11108 => y_in <= "10101011"; x_in <= "11100100"; z_correct<="0000100101001100";
        when 11109 => y_in <= "10101011"; x_in <= "11100101"; z_correct<="0000100011110111";
        when 11110 => y_in <= "10101011"; x_in <= "11100110"; z_correct<="0000100010100010";
        when 11111 => y_in <= "10101011"; x_in <= "11100111"; z_correct<="0000100001001101";
        when 11112 => y_in <= "10101011"; x_in <= "11101000"; z_correct<="0000011111111000";
        when 11113 => y_in <= "10101011"; x_in <= "11101001"; z_correct<="0000011110100011";
        when 11114 => y_in <= "10101011"; x_in <= "11101010"; z_correct<="0000011101001110";
        when 11115 => y_in <= "10101011"; x_in <= "11101011"; z_correct<="0000011011111001";
        when 11116 => y_in <= "10101011"; x_in <= "11101100"; z_correct<="0000011010100100";
        when 11117 => y_in <= "10101011"; x_in <= "11101101"; z_correct<="0000011001001111";
        when 11118 => y_in <= "10101011"; x_in <= "11101110"; z_correct<="0000010111111010";
        when 11119 => y_in <= "10101011"; x_in <= "11101111"; z_correct<="0000010110100101";
        when 11120 => y_in <= "10101011"; x_in <= "11110000"; z_correct<="0000010101010000";
        when 11121 => y_in <= "10101011"; x_in <= "11110001"; z_correct<="0000010011111011";
        when 11122 => y_in <= "10101011"; x_in <= "11110010"; z_correct<="0000010010100110";
        when 11123 => y_in <= "10101011"; x_in <= "11110011"; z_correct<="0000010001010001";
        when 11124 => y_in <= "10101011"; x_in <= "11110100"; z_correct<="0000001111111100";
        when 11125 => y_in <= "10101011"; x_in <= "11110101"; z_correct<="0000001110100111";
        when 11126 => y_in <= "10101011"; x_in <= "11110110"; z_correct<="0000001101010010";
        when 11127 => y_in <= "10101011"; x_in <= "11110111"; z_correct<="0000001011111101";
        when 11128 => y_in <= "10101011"; x_in <= "11111000"; z_correct<="0000001010101000";
        when 11129 => y_in <= "10101011"; x_in <= "11111001"; z_correct<="0000001001010011";
        when 11130 => y_in <= "10101011"; x_in <= "11111010"; z_correct<="0000000111111110";
        when 11131 => y_in <= "10101011"; x_in <= "11111011"; z_correct<="0000000110101001";
        when 11132 => y_in <= "10101011"; x_in <= "11111100"; z_correct<="0000000101010100";
        when 11133 => y_in <= "10101011"; x_in <= "11111101"; z_correct<="0000000011111111";
        when 11134 => y_in <= "10101011"; x_in <= "11111110"; z_correct<="0000000010101010";
        when 11135 => y_in <= "10101011"; x_in <= "11111111"; z_correct<="0000000001010101";
        when 11136 => y_in <= "10101011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 11137 => y_in <= "10101011"; x_in <= "00000001"; z_correct<="1111111110101011";
        when 11138 => y_in <= "10101011"; x_in <= "00000010"; z_correct<="1111111101010110";
        when 11139 => y_in <= "10101011"; x_in <= "00000011"; z_correct<="1111111100000001";
        when 11140 => y_in <= "10101011"; x_in <= "00000100"; z_correct<="1111111010101100";
        when 11141 => y_in <= "10101011"; x_in <= "00000101"; z_correct<="1111111001010111";
        when 11142 => y_in <= "10101011"; x_in <= "00000110"; z_correct<="1111111000000010";
        when 11143 => y_in <= "10101011"; x_in <= "00000111"; z_correct<="1111110110101101";
        when 11144 => y_in <= "10101011"; x_in <= "00001000"; z_correct<="1111110101011000";
        when 11145 => y_in <= "10101011"; x_in <= "00001001"; z_correct<="1111110100000011";
        when 11146 => y_in <= "10101011"; x_in <= "00001010"; z_correct<="1111110010101110";
        when 11147 => y_in <= "10101011"; x_in <= "00001011"; z_correct<="1111110001011001";
        when 11148 => y_in <= "10101011"; x_in <= "00001100"; z_correct<="1111110000000100";
        when 11149 => y_in <= "10101011"; x_in <= "00001101"; z_correct<="1111101110101111";
        when 11150 => y_in <= "10101011"; x_in <= "00001110"; z_correct<="1111101101011010";
        when 11151 => y_in <= "10101011"; x_in <= "00001111"; z_correct<="1111101100000101";
        when 11152 => y_in <= "10101011"; x_in <= "00010000"; z_correct<="1111101010110000";
        when 11153 => y_in <= "10101011"; x_in <= "00010001"; z_correct<="1111101001011011";
        when 11154 => y_in <= "10101011"; x_in <= "00010010"; z_correct<="1111101000000110";
        when 11155 => y_in <= "10101011"; x_in <= "00010011"; z_correct<="1111100110110001";
        when 11156 => y_in <= "10101011"; x_in <= "00010100"; z_correct<="1111100101011100";
        when 11157 => y_in <= "10101011"; x_in <= "00010101"; z_correct<="1111100100000111";
        when 11158 => y_in <= "10101011"; x_in <= "00010110"; z_correct<="1111100010110010";
        when 11159 => y_in <= "10101011"; x_in <= "00010111"; z_correct<="1111100001011101";
        when 11160 => y_in <= "10101011"; x_in <= "00011000"; z_correct<="1111100000001000";
        when 11161 => y_in <= "10101011"; x_in <= "00011001"; z_correct<="1111011110110011";
        when 11162 => y_in <= "10101011"; x_in <= "00011010"; z_correct<="1111011101011110";
        when 11163 => y_in <= "10101011"; x_in <= "00011011"; z_correct<="1111011100001001";
        when 11164 => y_in <= "10101011"; x_in <= "00011100"; z_correct<="1111011010110100";
        when 11165 => y_in <= "10101011"; x_in <= "00011101"; z_correct<="1111011001011111";
        when 11166 => y_in <= "10101011"; x_in <= "00011110"; z_correct<="1111011000001010";
        when 11167 => y_in <= "10101011"; x_in <= "00011111"; z_correct<="1111010110110101";
        when 11168 => y_in <= "10101011"; x_in <= "00100000"; z_correct<="1111010101100000";
        when 11169 => y_in <= "10101011"; x_in <= "00100001"; z_correct<="1111010100001011";
        when 11170 => y_in <= "10101011"; x_in <= "00100010"; z_correct<="1111010010110110";
        when 11171 => y_in <= "10101011"; x_in <= "00100011"; z_correct<="1111010001100001";
        when 11172 => y_in <= "10101011"; x_in <= "00100100"; z_correct<="1111010000001100";
        when 11173 => y_in <= "10101011"; x_in <= "00100101"; z_correct<="1111001110110111";
        when 11174 => y_in <= "10101011"; x_in <= "00100110"; z_correct<="1111001101100010";
        when 11175 => y_in <= "10101011"; x_in <= "00100111"; z_correct<="1111001100001101";
        when 11176 => y_in <= "10101011"; x_in <= "00101000"; z_correct<="1111001010111000";
        when 11177 => y_in <= "10101011"; x_in <= "00101001"; z_correct<="1111001001100011";
        when 11178 => y_in <= "10101011"; x_in <= "00101010"; z_correct<="1111001000001110";
        when 11179 => y_in <= "10101011"; x_in <= "00101011"; z_correct<="1111000110111001";
        when 11180 => y_in <= "10101011"; x_in <= "00101100"; z_correct<="1111000101100100";
        when 11181 => y_in <= "10101011"; x_in <= "00101101"; z_correct<="1111000100001111";
        when 11182 => y_in <= "10101011"; x_in <= "00101110"; z_correct<="1111000010111010";
        when 11183 => y_in <= "10101011"; x_in <= "00101111"; z_correct<="1111000001100101";
        when 11184 => y_in <= "10101011"; x_in <= "00110000"; z_correct<="1111000000010000";
        when 11185 => y_in <= "10101011"; x_in <= "00110001"; z_correct<="1110111110111011";
        when 11186 => y_in <= "10101011"; x_in <= "00110010"; z_correct<="1110111101100110";
        when 11187 => y_in <= "10101011"; x_in <= "00110011"; z_correct<="1110111100010001";
        when 11188 => y_in <= "10101011"; x_in <= "00110100"; z_correct<="1110111010111100";
        when 11189 => y_in <= "10101011"; x_in <= "00110101"; z_correct<="1110111001100111";
        when 11190 => y_in <= "10101011"; x_in <= "00110110"; z_correct<="1110111000010010";
        when 11191 => y_in <= "10101011"; x_in <= "00110111"; z_correct<="1110110110111101";
        when 11192 => y_in <= "10101011"; x_in <= "00111000"; z_correct<="1110110101101000";
        when 11193 => y_in <= "10101011"; x_in <= "00111001"; z_correct<="1110110100010011";
        when 11194 => y_in <= "10101011"; x_in <= "00111010"; z_correct<="1110110010111110";
        when 11195 => y_in <= "10101011"; x_in <= "00111011"; z_correct<="1110110001101001";
        when 11196 => y_in <= "10101011"; x_in <= "00111100"; z_correct<="1110110000010100";
        when 11197 => y_in <= "10101011"; x_in <= "00111101"; z_correct<="1110101110111111";
        when 11198 => y_in <= "10101011"; x_in <= "00111110"; z_correct<="1110101101101010";
        when 11199 => y_in <= "10101011"; x_in <= "00111111"; z_correct<="1110101100010101";
        when 11200 => y_in <= "10101011"; x_in <= "01000000"; z_correct<="1110101011000000";
        when 11201 => y_in <= "10101011"; x_in <= "01000001"; z_correct<="1110101001101011";
        when 11202 => y_in <= "10101011"; x_in <= "01000010"; z_correct<="1110101000010110";
        when 11203 => y_in <= "10101011"; x_in <= "01000011"; z_correct<="1110100111000001";
        when 11204 => y_in <= "10101011"; x_in <= "01000100"; z_correct<="1110100101101100";
        when 11205 => y_in <= "10101011"; x_in <= "01000101"; z_correct<="1110100100010111";
        when 11206 => y_in <= "10101011"; x_in <= "01000110"; z_correct<="1110100011000010";
        when 11207 => y_in <= "10101011"; x_in <= "01000111"; z_correct<="1110100001101101";
        when 11208 => y_in <= "10101011"; x_in <= "01001000"; z_correct<="1110100000011000";
        when 11209 => y_in <= "10101011"; x_in <= "01001001"; z_correct<="1110011111000011";
        when 11210 => y_in <= "10101011"; x_in <= "01001010"; z_correct<="1110011101101110";
        when 11211 => y_in <= "10101011"; x_in <= "01001011"; z_correct<="1110011100011001";
        when 11212 => y_in <= "10101011"; x_in <= "01001100"; z_correct<="1110011011000100";
        when 11213 => y_in <= "10101011"; x_in <= "01001101"; z_correct<="1110011001101111";
        when 11214 => y_in <= "10101011"; x_in <= "01001110"; z_correct<="1110011000011010";
        when 11215 => y_in <= "10101011"; x_in <= "01001111"; z_correct<="1110010111000101";
        when 11216 => y_in <= "10101011"; x_in <= "01010000"; z_correct<="1110010101110000";
        when 11217 => y_in <= "10101011"; x_in <= "01010001"; z_correct<="1110010100011011";
        when 11218 => y_in <= "10101011"; x_in <= "01010010"; z_correct<="1110010011000110";
        when 11219 => y_in <= "10101011"; x_in <= "01010011"; z_correct<="1110010001110001";
        when 11220 => y_in <= "10101011"; x_in <= "01010100"; z_correct<="1110010000011100";
        when 11221 => y_in <= "10101011"; x_in <= "01010101"; z_correct<="1110001111000111";
        when 11222 => y_in <= "10101011"; x_in <= "01010110"; z_correct<="1110001101110010";
        when 11223 => y_in <= "10101011"; x_in <= "01010111"; z_correct<="1110001100011101";
        when 11224 => y_in <= "10101011"; x_in <= "01011000"; z_correct<="1110001011001000";
        when 11225 => y_in <= "10101011"; x_in <= "01011001"; z_correct<="1110001001110011";
        when 11226 => y_in <= "10101011"; x_in <= "01011010"; z_correct<="1110001000011110";
        when 11227 => y_in <= "10101011"; x_in <= "01011011"; z_correct<="1110000111001001";
        when 11228 => y_in <= "10101011"; x_in <= "01011100"; z_correct<="1110000101110100";
        when 11229 => y_in <= "10101011"; x_in <= "01011101"; z_correct<="1110000100011111";
        when 11230 => y_in <= "10101011"; x_in <= "01011110"; z_correct<="1110000011001010";
        when 11231 => y_in <= "10101011"; x_in <= "01011111"; z_correct<="1110000001110101";
        when 11232 => y_in <= "10101011"; x_in <= "01100000"; z_correct<="1110000000100000";
        when 11233 => y_in <= "10101011"; x_in <= "01100001"; z_correct<="1101111111001011";
        when 11234 => y_in <= "10101011"; x_in <= "01100010"; z_correct<="1101111101110110";
        when 11235 => y_in <= "10101011"; x_in <= "01100011"; z_correct<="1101111100100001";
        when 11236 => y_in <= "10101011"; x_in <= "01100100"; z_correct<="1101111011001100";
        when 11237 => y_in <= "10101011"; x_in <= "01100101"; z_correct<="1101111001110111";
        when 11238 => y_in <= "10101011"; x_in <= "01100110"; z_correct<="1101111000100010";
        when 11239 => y_in <= "10101011"; x_in <= "01100111"; z_correct<="1101110111001101";
        when 11240 => y_in <= "10101011"; x_in <= "01101000"; z_correct<="1101110101111000";
        when 11241 => y_in <= "10101011"; x_in <= "01101001"; z_correct<="1101110100100011";
        when 11242 => y_in <= "10101011"; x_in <= "01101010"; z_correct<="1101110011001110";
        when 11243 => y_in <= "10101011"; x_in <= "01101011"; z_correct<="1101110001111001";
        when 11244 => y_in <= "10101011"; x_in <= "01101100"; z_correct<="1101110000100100";
        when 11245 => y_in <= "10101011"; x_in <= "01101101"; z_correct<="1101101111001111";
        when 11246 => y_in <= "10101011"; x_in <= "01101110"; z_correct<="1101101101111010";
        when 11247 => y_in <= "10101011"; x_in <= "01101111"; z_correct<="1101101100100101";
        when 11248 => y_in <= "10101011"; x_in <= "01110000"; z_correct<="1101101011010000";
        when 11249 => y_in <= "10101011"; x_in <= "01110001"; z_correct<="1101101001111011";
        when 11250 => y_in <= "10101011"; x_in <= "01110010"; z_correct<="1101101000100110";
        when 11251 => y_in <= "10101011"; x_in <= "01110011"; z_correct<="1101100111010001";
        when 11252 => y_in <= "10101011"; x_in <= "01110100"; z_correct<="1101100101111100";
        when 11253 => y_in <= "10101011"; x_in <= "01110101"; z_correct<="1101100100100111";
        when 11254 => y_in <= "10101011"; x_in <= "01110110"; z_correct<="1101100011010010";
        when 11255 => y_in <= "10101011"; x_in <= "01110111"; z_correct<="1101100001111101";
        when 11256 => y_in <= "10101011"; x_in <= "01111000"; z_correct<="1101100000101000";
        when 11257 => y_in <= "10101011"; x_in <= "01111001"; z_correct<="1101011111010011";
        when 11258 => y_in <= "10101011"; x_in <= "01111010"; z_correct<="1101011101111110";
        when 11259 => y_in <= "10101011"; x_in <= "01111011"; z_correct<="1101011100101001";
        when 11260 => y_in <= "10101011"; x_in <= "01111100"; z_correct<="1101011011010100";
        when 11261 => y_in <= "10101011"; x_in <= "01111101"; z_correct<="1101011001111111";
        when 11262 => y_in <= "10101011"; x_in <= "01111110"; z_correct<="1101011000101010";
        when 11263 => y_in <= "10101011"; x_in <= "01111111"; z_correct<="1101010111010101";
        when 11264 => y_in <= "10101100"; x_in <= "10000000"; z_correct<="0010101000000000";
        when 11265 => y_in <= "10101100"; x_in <= "10000001"; z_correct<="0010100110101100";
        when 11266 => y_in <= "10101100"; x_in <= "10000010"; z_correct<="0010100101011000";
        when 11267 => y_in <= "10101100"; x_in <= "10000011"; z_correct<="0010100100000100";
        when 11268 => y_in <= "10101100"; x_in <= "10000100"; z_correct<="0010100010110000";
        when 11269 => y_in <= "10101100"; x_in <= "10000101"; z_correct<="0010100001011100";
        when 11270 => y_in <= "10101100"; x_in <= "10000110"; z_correct<="0010100000001000";
        when 11271 => y_in <= "10101100"; x_in <= "10000111"; z_correct<="0010011110110100";
        when 11272 => y_in <= "10101100"; x_in <= "10001000"; z_correct<="0010011101100000";
        when 11273 => y_in <= "10101100"; x_in <= "10001001"; z_correct<="0010011100001100";
        when 11274 => y_in <= "10101100"; x_in <= "10001010"; z_correct<="0010011010111000";
        when 11275 => y_in <= "10101100"; x_in <= "10001011"; z_correct<="0010011001100100";
        when 11276 => y_in <= "10101100"; x_in <= "10001100"; z_correct<="0010011000010000";
        when 11277 => y_in <= "10101100"; x_in <= "10001101"; z_correct<="0010010110111100";
        when 11278 => y_in <= "10101100"; x_in <= "10001110"; z_correct<="0010010101101000";
        when 11279 => y_in <= "10101100"; x_in <= "10001111"; z_correct<="0010010100010100";
        when 11280 => y_in <= "10101100"; x_in <= "10010000"; z_correct<="0010010011000000";
        when 11281 => y_in <= "10101100"; x_in <= "10010001"; z_correct<="0010010001101100";
        when 11282 => y_in <= "10101100"; x_in <= "10010010"; z_correct<="0010010000011000";
        when 11283 => y_in <= "10101100"; x_in <= "10010011"; z_correct<="0010001111000100";
        when 11284 => y_in <= "10101100"; x_in <= "10010100"; z_correct<="0010001101110000";
        when 11285 => y_in <= "10101100"; x_in <= "10010101"; z_correct<="0010001100011100";
        when 11286 => y_in <= "10101100"; x_in <= "10010110"; z_correct<="0010001011001000";
        when 11287 => y_in <= "10101100"; x_in <= "10010111"; z_correct<="0010001001110100";
        when 11288 => y_in <= "10101100"; x_in <= "10011000"; z_correct<="0010001000100000";
        when 11289 => y_in <= "10101100"; x_in <= "10011001"; z_correct<="0010000111001100";
        when 11290 => y_in <= "10101100"; x_in <= "10011010"; z_correct<="0010000101111000";
        when 11291 => y_in <= "10101100"; x_in <= "10011011"; z_correct<="0010000100100100";
        when 11292 => y_in <= "10101100"; x_in <= "10011100"; z_correct<="0010000011010000";
        when 11293 => y_in <= "10101100"; x_in <= "10011101"; z_correct<="0010000001111100";
        when 11294 => y_in <= "10101100"; x_in <= "10011110"; z_correct<="0010000000101000";
        when 11295 => y_in <= "10101100"; x_in <= "10011111"; z_correct<="0001111111010100";
        when 11296 => y_in <= "10101100"; x_in <= "10100000"; z_correct<="0001111110000000";
        when 11297 => y_in <= "10101100"; x_in <= "10100001"; z_correct<="0001111100101100";
        when 11298 => y_in <= "10101100"; x_in <= "10100010"; z_correct<="0001111011011000";
        when 11299 => y_in <= "10101100"; x_in <= "10100011"; z_correct<="0001111010000100";
        when 11300 => y_in <= "10101100"; x_in <= "10100100"; z_correct<="0001111000110000";
        when 11301 => y_in <= "10101100"; x_in <= "10100101"; z_correct<="0001110111011100";
        when 11302 => y_in <= "10101100"; x_in <= "10100110"; z_correct<="0001110110001000";
        when 11303 => y_in <= "10101100"; x_in <= "10100111"; z_correct<="0001110100110100";
        when 11304 => y_in <= "10101100"; x_in <= "10101000"; z_correct<="0001110011100000";
        when 11305 => y_in <= "10101100"; x_in <= "10101001"; z_correct<="0001110010001100";
        when 11306 => y_in <= "10101100"; x_in <= "10101010"; z_correct<="0001110000111000";
        when 11307 => y_in <= "10101100"; x_in <= "10101011"; z_correct<="0001101111100100";
        when 11308 => y_in <= "10101100"; x_in <= "10101100"; z_correct<="0001101110010000";
        when 11309 => y_in <= "10101100"; x_in <= "10101101"; z_correct<="0001101100111100";
        when 11310 => y_in <= "10101100"; x_in <= "10101110"; z_correct<="0001101011101000";
        when 11311 => y_in <= "10101100"; x_in <= "10101111"; z_correct<="0001101010010100";
        when 11312 => y_in <= "10101100"; x_in <= "10110000"; z_correct<="0001101001000000";
        when 11313 => y_in <= "10101100"; x_in <= "10110001"; z_correct<="0001100111101100";
        when 11314 => y_in <= "10101100"; x_in <= "10110010"; z_correct<="0001100110011000";
        when 11315 => y_in <= "10101100"; x_in <= "10110011"; z_correct<="0001100101000100";
        when 11316 => y_in <= "10101100"; x_in <= "10110100"; z_correct<="0001100011110000";
        when 11317 => y_in <= "10101100"; x_in <= "10110101"; z_correct<="0001100010011100";
        when 11318 => y_in <= "10101100"; x_in <= "10110110"; z_correct<="0001100001001000";
        when 11319 => y_in <= "10101100"; x_in <= "10110111"; z_correct<="0001011111110100";
        when 11320 => y_in <= "10101100"; x_in <= "10111000"; z_correct<="0001011110100000";
        when 11321 => y_in <= "10101100"; x_in <= "10111001"; z_correct<="0001011101001100";
        when 11322 => y_in <= "10101100"; x_in <= "10111010"; z_correct<="0001011011111000";
        when 11323 => y_in <= "10101100"; x_in <= "10111011"; z_correct<="0001011010100100";
        when 11324 => y_in <= "10101100"; x_in <= "10111100"; z_correct<="0001011001010000";
        when 11325 => y_in <= "10101100"; x_in <= "10111101"; z_correct<="0001010111111100";
        when 11326 => y_in <= "10101100"; x_in <= "10111110"; z_correct<="0001010110101000";
        when 11327 => y_in <= "10101100"; x_in <= "10111111"; z_correct<="0001010101010100";
        when 11328 => y_in <= "10101100"; x_in <= "11000000"; z_correct<="0001010100000000";
        when 11329 => y_in <= "10101100"; x_in <= "11000001"; z_correct<="0001010010101100";
        when 11330 => y_in <= "10101100"; x_in <= "11000010"; z_correct<="0001010001011000";
        when 11331 => y_in <= "10101100"; x_in <= "11000011"; z_correct<="0001010000000100";
        when 11332 => y_in <= "10101100"; x_in <= "11000100"; z_correct<="0001001110110000";
        when 11333 => y_in <= "10101100"; x_in <= "11000101"; z_correct<="0001001101011100";
        when 11334 => y_in <= "10101100"; x_in <= "11000110"; z_correct<="0001001100001000";
        when 11335 => y_in <= "10101100"; x_in <= "11000111"; z_correct<="0001001010110100";
        when 11336 => y_in <= "10101100"; x_in <= "11001000"; z_correct<="0001001001100000";
        when 11337 => y_in <= "10101100"; x_in <= "11001001"; z_correct<="0001001000001100";
        when 11338 => y_in <= "10101100"; x_in <= "11001010"; z_correct<="0001000110111000";
        when 11339 => y_in <= "10101100"; x_in <= "11001011"; z_correct<="0001000101100100";
        when 11340 => y_in <= "10101100"; x_in <= "11001100"; z_correct<="0001000100010000";
        when 11341 => y_in <= "10101100"; x_in <= "11001101"; z_correct<="0001000010111100";
        when 11342 => y_in <= "10101100"; x_in <= "11001110"; z_correct<="0001000001101000";
        when 11343 => y_in <= "10101100"; x_in <= "11001111"; z_correct<="0001000000010100";
        when 11344 => y_in <= "10101100"; x_in <= "11010000"; z_correct<="0000111111000000";
        when 11345 => y_in <= "10101100"; x_in <= "11010001"; z_correct<="0000111101101100";
        when 11346 => y_in <= "10101100"; x_in <= "11010010"; z_correct<="0000111100011000";
        when 11347 => y_in <= "10101100"; x_in <= "11010011"; z_correct<="0000111011000100";
        when 11348 => y_in <= "10101100"; x_in <= "11010100"; z_correct<="0000111001110000";
        when 11349 => y_in <= "10101100"; x_in <= "11010101"; z_correct<="0000111000011100";
        when 11350 => y_in <= "10101100"; x_in <= "11010110"; z_correct<="0000110111001000";
        when 11351 => y_in <= "10101100"; x_in <= "11010111"; z_correct<="0000110101110100";
        when 11352 => y_in <= "10101100"; x_in <= "11011000"; z_correct<="0000110100100000";
        when 11353 => y_in <= "10101100"; x_in <= "11011001"; z_correct<="0000110011001100";
        when 11354 => y_in <= "10101100"; x_in <= "11011010"; z_correct<="0000110001111000";
        when 11355 => y_in <= "10101100"; x_in <= "11011011"; z_correct<="0000110000100100";
        when 11356 => y_in <= "10101100"; x_in <= "11011100"; z_correct<="0000101111010000";
        when 11357 => y_in <= "10101100"; x_in <= "11011101"; z_correct<="0000101101111100";
        when 11358 => y_in <= "10101100"; x_in <= "11011110"; z_correct<="0000101100101000";
        when 11359 => y_in <= "10101100"; x_in <= "11011111"; z_correct<="0000101011010100";
        when 11360 => y_in <= "10101100"; x_in <= "11100000"; z_correct<="0000101010000000";
        when 11361 => y_in <= "10101100"; x_in <= "11100001"; z_correct<="0000101000101100";
        when 11362 => y_in <= "10101100"; x_in <= "11100010"; z_correct<="0000100111011000";
        when 11363 => y_in <= "10101100"; x_in <= "11100011"; z_correct<="0000100110000100";
        when 11364 => y_in <= "10101100"; x_in <= "11100100"; z_correct<="0000100100110000";
        when 11365 => y_in <= "10101100"; x_in <= "11100101"; z_correct<="0000100011011100";
        when 11366 => y_in <= "10101100"; x_in <= "11100110"; z_correct<="0000100010001000";
        when 11367 => y_in <= "10101100"; x_in <= "11100111"; z_correct<="0000100000110100";
        when 11368 => y_in <= "10101100"; x_in <= "11101000"; z_correct<="0000011111100000";
        when 11369 => y_in <= "10101100"; x_in <= "11101001"; z_correct<="0000011110001100";
        when 11370 => y_in <= "10101100"; x_in <= "11101010"; z_correct<="0000011100111000";
        when 11371 => y_in <= "10101100"; x_in <= "11101011"; z_correct<="0000011011100100";
        when 11372 => y_in <= "10101100"; x_in <= "11101100"; z_correct<="0000011010010000";
        when 11373 => y_in <= "10101100"; x_in <= "11101101"; z_correct<="0000011000111100";
        when 11374 => y_in <= "10101100"; x_in <= "11101110"; z_correct<="0000010111101000";
        when 11375 => y_in <= "10101100"; x_in <= "11101111"; z_correct<="0000010110010100";
        when 11376 => y_in <= "10101100"; x_in <= "11110000"; z_correct<="0000010101000000";
        when 11377 => y_in <= "10101100"; x_in <= "11110001"; z_correct<="0000010011101100";
        when 11378 => y_in <= "10101100"; x_in <= "11110010"; z_correct<="0000010010011000";
        when 11379 => y_in <= "10101100"; x_in <= "11110011"; z_correct<="0000010001000100";
        when 11380 => y_in <= "10101100"; x_in <= "11110100"; z_correct<="0000001111110000";
        when 11381 => y_in <= "10101100"; x_in <= "11110101"; z_correct<="0000001110011100";
        when 11382 => y_in <= "10101100"; x_in <= "11110110"; z_correct<="0000001101001000";
        when 11383 => y_in <= "10101100"; x_in <= "11110111"; z_correct<="0000001011110100";
        when 11384 => y_in <= "10101100"; x_in <= "11111000"; z_correct<="0000001010100000";
        when 11385 => y_in <= "10101100"; x_in <= "11111001"; z_correct<="0000001001001100";
        when 11386 => y_in <= "10101100"; x_in <= "11111010"; z_correct<="0000000111111000";
        when 11387 => y_in <= "10101100"; x_in <= "11111011"; z_correct<="0000000110100100";
        when 11388 => y_in <= "10101100"; x_in <= "11111100"; z_correct<="0000000101010000";
        when 11389 => y_in <= "10101100"; x_in <= "11111101"; z_correct<="0000000011111100";
        when 11390 => y_in <= "10101100"; x_in <= "11111110"; z_correct<="0000000010101000";
        when 11391 => y_in <= "10101100"; x_in <= "11111111"; z_correct<="0000000001010100";
        when 11392 => y_in <= "10101100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 11393 => y_in <= "10101100"; x_in <= "00000001"; z_correct<="1111111110101100";
        when 11394 => y_in <= "10101100"; x_in <= "00000010"; z_correct<="1111111101011000";
        when 11395 => y_in <= "10101100"; x_in <= "00000011"; z_correct<="1111111100000100";
        when 11396 => y_in <= "10101100"; x_in <= "00000100"; z_correct<="1111111010110000";
        when 11397 => y_in <= "10101100"; x_in <= "00000101"; z_correct<="1111111001011100";
        when 11398 => y_in <= "10101100"; x_in <= "00000110"; z_correct<="1111111000001000";
        when 11399 => y_in <= "10101100"; x_in <= "00000111"; z_correct<="1111110110110100";
        when 11400 => y_in <= "10101100"; x_in <= "00001000"; z_correct<="1111110101100000";
        when 11401 => y_in <= "10101100"; x_in <= "00001001"; z_correct<="1111110100001100";
        when 11402 => y_in <= "10101100"; x_in <= "00001010"; z_correct<="1111110010111000";
        when 11403 => y_in <= "10101100"; x_in <= "00001011"; z_correct<="1111110001100100";
        when 11404 => y_in <= "10101100"; x_in <= "00001100"; z_correct<="1111110000010000";
        when 11405 => y_in <= "10101100"; x_in <= "00001101"; z_correct<="1111101110111100";
        when 11406 => y_in <= "10101100"; x_in <= "00001110"; z_correct<="1111101101101000";
        when 11407 => y_in <= "10101100"; x_in <= "00001111"; z_correct<="1111101100010100";
        when 11408 => y_in <= "10101100"; x_in <= "00010000"; z_correct<="1111101011000000";
        when 11409 => y_in <= "10101100"; x_in <= "00010001"; z_correct<="1111101001101100";
        when 11410 => y_in <= "10101100"; x_in <= "00010010"; z_correct<="1111101000011000";
        when 11411 => y_in <= "10101100"; x_in <= "00010011"; z_correct<="1111100111000100";
        when 11412 => y_in <= "10101100"; x_in <= "00010100"; z_correct<="1111100101110000";
        when 11413 => y_in <= "10101100"; x_in <= "00010101"; z_correct<="1111100100011100";
        when 11414 => y_in <= "10101100"; x_in <= "00010110"; z_correct<="1111100011001000";
        when 11415 => y_in <= "10101100"; x_in <= "00010111"; z_correct<="1111100001110100";
        when 11416 => y_in <= "10101100"; x_in <= "00011000"; z_correct<="1111100000100000";
        when 11417 => y_in <= "10101100"; x_in <= "00011001"; z_correct<="1111011111001100";
        when 11418 => y_in <= "10101100"; x_in <= "00011010"; z_correct<="1111011101111000";
        when 11419 => y_in <= "10101100"; x_in <= "00011011"; z_correct<="1111011100100100";
        when 11420 => y_in <= "10101100"; x_in <= "00011100"; z_correct<="1111011011010000";
        when 11421 => y_in <= "10101100"; x_in <= "00011101"; z_correct<="1111011001111100";
        when 11422 => y_in <= "10101100"; x_in <= "00011110"; z_correct<="1111011000101000";
        when 11423 => y_in <= "10101100"; x_in <= "00011111"; z_correct<="1111010111010100";
        when 11424 => y_in <= "10101100"; x_in <= "00100000"; z_correct<="1111010110000000";
        when 11425 => y_in <= "10101100"; x_in <= "00100001"; z_correct<="1111010100101100";
        when 11426 => y_in <= "10101100"; x_in <= "00100010"; z_correct<="1111010011011000";
        when 11427 => y_in <= "10101100"; x_in <= "00100011"; z_correct<="1111010010000100";
        when 11428 => y_in <= "10101100"; x_in <= "00100100"; z_correct<="1111010000110000";
        when 11429 => y_in <= "10101100"; x_in <= "00100101"; z_correct<="1111001111011100";
        when 11430 => y_in <= "10101100"; x_in <= "00100110"; z_correct<="1111001110001000";
        when 11431 => y_in <= "10101100"; x_in <= "00100111"; z_correct<="1111001100110100";
        when 11432 => y_in <= "10101100"; x_in <= "00101000"; z_correct<="1111001011100000";
        when 11433 => y_in <= "10101100"; x_in <= "00101001"; z_correct<="1111001010001100";
        when 11434 => y_in <= "10101100"; x_in <= "00101010"; z_correct<="1111001000111000";
        when 11435 => y_in <= "10101100"; x_in <= "00101011"; z_correct<="1111000111100100";
        when 11436 => y_in <= "10101100"; x_in <= "00101100"; z_correct<="1111000110010000";
        when 11437 => y_in <= "10101100"; x_in <= "00101101"; z_correct<="1111000100111100";
        when 11438 => y_in <= "10101100"; x_in <= "00101110"; z_correct<="1111000011101000";
        when 11439 => y_in <= "10101100"; x_in <= "00101111"; z_correct<="1111000010010100";
        when 11440 => y_in <= "10101100"; x_in <= "00110000"; z_correct<="1111000001000000";
        when 11441 => y_in <= "10101100"; x_in <= "00110001"; z_correct<="1110111111101100";
        when 11442 => y_in <= "10101100"; x_in <= "00110010"; z_correct<="1110111110011000";
        when 11443 => y_in <= "10101100"; x_in <= "00110011"; z_correct<="1110111101000100";
        when 11444 => y_in <= "10101100"; x_in <= "00110100"; z_correct<="1110111011110000";
        when 11445 => y_in <= "10101100"; x_in <= "00110101"; z_correct<="1110111010011100";
        when 11446 => y_in <= "10101100"; x_in <= "00110110"; z_correct<="1110111001001000";
        when 11447 => y_in <= "10101100"; x_in <= "00110111"; z_correct<="1110110111110100";
        when 11448 => y_in <= "10101100"; x_in <= "00111000"; z_correct<="1110110110100000";
        when 11449 => y_in <= "10101100"; x_in <= "00111001"; z_correct<="1110110101001100";
        when 11450 => y_in <= "10101100"; x_in <= "00111010"; z_correct<="1110110011111000";
        when 11451 => y_in <= "10101100"; x_in <= "00111011"; z_correct<="1110110010100100";
        when 11452 => y_in <= "10101100"; x_in <= "00111100"; z_correct<="1110110001010000";
        when 11453 => y_in <= "10101100"; x_in <= "00111101"; z_correct<="1110101111111100";
        when 11454 => y_in <= "10101100"; x_in <= "00111110"; z_correct<="1110101110101000";
        when 11455 => y_in <= "10101100"; x_in <= "00111111"; z_correct<="1110101101010100";
        when 11456 => y_in <= "10101100"; x_in <= "01000000"; z_correct<="1110101100000000";
        when 11457 => y_in <= "10101100"; x_in <= "01000001"; z_correct<="1110101010101100";
        when 11458 => y_in <= "10101100"; x_in <= "01000010"; z_correct<="1110101001011000";
        when 11459 => y_in <= "10101100"; x_in <= "01000011"; z_correct<="1110101000000100";
        when 11460 => y_in <= "10101100"; x_in <= "01000100"; z_correct<="1110100110110000";
        when 11461 => y_in <= "10101100"; x_in <= "01000101"; z_correct<="1110100101011100";
        when 11462 => y_in <= "10101100"; x_in <= "01000110"; z_correct<="1110100100001000";
        when 11463 => y_in <= "10101100"; x_in <= "01000111"; z_correct<="1110100010110100";
        when 11464 => y_in <= "10101100"; x_in <= "01001000"; z_correct<="1110100001100000";
        when 11465 => y_in <= "10101100"; x_in <= "01001001"; z_correct<="1110100000001100";
        when 11466 => y_in <= "10101100"; x_in <= "01001010"; z_correct<="1110011110111000";
        when 11467 => y_in <= "10101100"; x_in <= "01001011"; z_correct<="1110011101100100";
        when 11468 => y_in <= "10101100"; x_in <= "01001100"; z_correct<="1110011100010000";
        when 11469 => y_in <= "10101100"; x_in <= "01001101"; z_correct<="1110011010111100";
        when 11470 => y_in <= "10101100"; x_in <= "01001110"; z_correct<="1110011001101000";
        when 11471 => y_in <= "10101100"; x_in <= "01001111"; z_correct<="1110011000010100";
        when 11472 => y_in <= "10101100"; x_in <= "01010000"; z_correct<="1110010111000000";
        when 11473 => y_in <= "10101100"; x_in <= "01010001"; z_correct<="1110010101101100";
        when 11474 => y_in <= "10101100"; x_in <= "01010010"; z_correct<="1110010100011000";
        when 11475 => y_in <= "10101100"; x_in <= "01010011"; z_correct<="1110010011000100";
        when 11476 => y_in <= "10101100"; x_in <= "01010100"; z_correct<="1110010001110000";
        when 11477 => y_in <= "10101100"; x_in <= "01010101"; z_correct<="1110010000011100";
        when 11478 => y_in <= "10101100"; x_in <= "01010110"; z_correct<="1110001111001000";
        when 11479 => y_in <= "10101100"; x_in <= "01010111"; z_correct<="1110001101110100";
        when 11480 => y_in <= "10101100"; x_in <= "01011000"; z_correct<="1110001100100000";
        when 11481 => y_in <= "10101100"; x_in <= "01011001"; z_correct<="1110001011001100";
        when 11482 => y_in <= "10101100"; x_in <= "01011010"; z_correct<="1110001001111000";
        when 11483 => y_in <= "10101100"; x_in <= "01011011"; z_correct<="1110001000100100";
        when 11484 => y_in <= "10101100"; x_in <= "01011100"; z_correct<="1110000111010000";
        when 11485 => y_in <= "10101100"; x_in <= "01011101"; z_correct<="1110000101111100";
        when 11486 => y_in <= "10101100"; x_in <= "01011110"; z_correct<="1110000100101000";
        when 11487 => y_in <= "10101100"; x_in <= "01011111"; z_correct<="1110000011010100";
        when 11488 => y_in <= "10101100"; x_in <= "01100000"; z_correct<="1110000010000000";
        when 11489 => y_in <= "10101100"; x_in <= "01100001"; z_correct<="1110000000101100";
        when 11490 => y_in <= "10101100"; x_in <= "01100010"; z_correct<="1101111111011000";
        when 11491 => y_in <= "10101100"; x_in <= "01100011"; z_correct<="1101111110000100";
        when 11492 => y_in <= "10101100"; x_in <= "01100100"; z_correct<="1101111100110000";
        when 11493 => y_in <= "10101100"; x_in <= "01100101"; z_correct<="1101111011011100";
        when 11494 => y_in <= "10101100"; x_in <= "01100110"; z_correct<="1101111010001000";
        when 11495 => y_in <= "10101100"; x_in <= "01100111"; z_correct<="1101111000110100";
        when 11496 => y_in <= "10101100"; x_in <= "01101000"; z_correct<="1101110111100000";
        when 11497 => y_in <= "10101100"; x_in <= "01101001"; z_correct<="1101110110001100";
        when 11498 => y_in <= "10101100"; x_in <= "01101010"; z_correct<="1101110100111000";
        when 11499 => y_in <= "10101100"; x_in <= "01101011"; z_correct<="1101110011100100";
        when 11500 => y_in <= "10101100"; x_in <= "01101100"; z_correct<="1101110010010000";
        when 11501 => y_in <= "10101100"; x_in <= "01101101"; z_correct<="1101110000111100";
        when 11502 => y_in <= "10101100"; x_in <= "01101110"; z_correct<="1101101111101000";
        when 11503 => y_in <= "10101100"; x_in <= "01101111"; z_correct<="1101101110010100";
        when 11504 => y_in <= "10101100"; x_in <= "01110000"; z_correct<="1101101101000000";
        when 11505 => y_in <= "10101100"; x_in <= "01110001"; z_correct<="1101101011101100";
        when 11506 => y_in <= "10101100"; x_in <= "01110010"; z_correct<="1101101010011000";
        when 11507 => y_in <= "10101100"; x_in <= "01110011"; z_correct<="1101101001000100";
        when 11508 => y_in <= "10101100"; x_in <= "01110100"; z_correct<="1101100111110000";
        when 11509 => y_in <= "10101100"; x_in <= "01110101"; z_correct<="1101100110011100";
        when 11510 => y_in <= "10101100"; x_in <= "01110110"; z_correct<="1101100101001000";
        when 11511 => y_in <= "10101100"; x_in <= "01110111"; z_correct<="1101100011110100";
        when 11512 => y_in <= "10101100"; x_in <= "01111000"; z_correct<="1101100010100000";
        when 11513 => y_in <= "10101100"; x_in <= "01111001"; z_correct<="1101100001001100";
        when 11514 => y_in <= "10101100"; x_in <= "01111010"; z_correct<="1101011111111000";
        when 11515 => y_in <= "10101100"; x_in <= "01111011"; z_correct<="1101011110100100";
        when 11516 => y_in <= "10101100"; x_in <= "01111100"; z_correct<="1101011101010000";
        when 11517 => y_in <= "10101100"; x_in <= "01111101"; z_correct<="1101011011111100";
        when 11518 => y_in <= "10101100"; x_in <= "01111110"; z_correct<="1101011010101000";
        when 11519 => y_in <= "10101100"; x_in <= "01111111"; z_correct<="1101011001010100";
        when 11520 => y_in <= "10101101"; x_in <= "10000000"; z_correct<="0010100110000000";
        when 11521 => y_in <= "10101101"; x_in <= "10000001"; z_correct<="0010100100101101";
        when 11522 => y_in <= "10101101"; x_in <= "10000010"; z_correct<="0010100011011010";
        when 11523 => y_in <= "10101101"; x_in <= "10000011"; z_correct<="0010100010000111";
        when 11524 => y_in <= "10101101"; x_in <= "10000100"; z_correct<="0010100000110100";
        when 11525 => y_in <= "10101101"; x_in <= "10000101"; z_correct<="0010011111100001";
        when 11526 => y_in <= "10101101"; x_in <= "10000110"; z_correct<="0010011110001110";
        when 11527 => y_in <= "10101101"; x_in <= "10000111"; z_correct<="0010011100111011";
        when 11528 => y_in <= "10101101"; x_in <= "10001000"; z_correct<="0010011011101000";
        when 11529 => y_in <= "10101101"; x_in <= "10001001"; z_correct<="0010011010010101";
        when 11530 => y_in <= "10101101"; x_in <= "10001010"; z_correct<="0010011001000010";
        when 11531 => y_in <= "10101101"; x_in <= "10001011"; z_correct<="0010010111101111";
        when 11532 => y_in <= "10101101"; x_in <= "10001100"; z_correct<="0010010110011100";
        when 11533 => y_in <= "10101101"; x_in <= "10001101"; z_correct<="0010010101001001";
        when 11534 => y_in <= "10101101"; x_in <= "10001110"; z_correct<="0010010011110110";
        when 11535 => y_in <= "10101101"; x_in <= "10001111"; z_correct<="0010010010100011";
        when 11536 => y_in <= "10101101"; x_in <= "10010000"; z_correct<="0010010001010000";
        when 11537 => y_in <= "10101101"; x_in <= "10010001"; z_correct<="0010001111111101";
        when 11538 => y_in <= "10101101"; x_in <= "10010010"; z_correct<="0010001110101010";
        when 11539 => y_in <= "10101101"; x_in <= "10010011"; z_correct<="0010001101010111";
        when 11540 => y_in <= "10101101"; x_in <= "10010100"; z_correct<="0010001100000100";
        when 11541 => y_in <= "10101101"; x_in <= "10010101"; z_correct<="0010001010110001";
        when 11542 => y_in <= "10101101"; x_in <= "10010110"; z_correct<="0010001001011110";
        when 11543 => y_in <= "10101101"; x_in <= "10010111"; z_correct<="0010001000001011";
        when 11544 => y_in <= "10101101"; x_in <= "10011000"; z_correct<="0010000110111000";
        when 11545 => y_in <= "10101101"; x_in <= "10011001"; z_correct<="0010000101100101";
        when 11546 => y_in <= "10101101"; x_in <= "10011010"; z_correct<="0010000100010010";
        when 11547 => y_in <= "10101101"; x_in <= "10011011"; z_correct<="0010000010111111";
        when 11548 => y_in <= "10101101"; x_in <= "10011100"; z_correct<="0010000001101100";
        when 11549 => y_in <= "10101101"; x_in <= "10011101"; z_correct<="0010000000011001";
        when 11550 => y_in <= "10101101"; x_in <= "10011110"; z_correct<="0001111111000110";
        when 11551 => y_in <= "10101101"; x_in <= "10011111"; z_correct<="0001111101110011";
        when 11552 => y_in <= "10101101"; x_in <= "10100000"; z_correct<="0001111100100000";
        when 11553 => y_in <= "10101101"; x_in <= "10100001"; z_correct<="0001111011001101";
        when 11554 => y_in <= "10101101"; x_in <= "10100010"; z_correct<="0001111001111010";
        when 11555 => y_in <= "10101101"; x_in <= "10100011"; z_correct<="0001111000100111";
        when 11556 => y_in <= "10101101"; x_in <= "10100100"; z_correct<="0001110111010100";
        when 11557 => y_in <= "10101101"; x_in <= "10100101"; z_correct<="0001110110000001";
        when 11558 => y_in <= "10101101"; x_in <= "10100110"; z_correct<="0001110100101110";
        when 11559 => y_in <= "10101101"; x_in <= "10100111"; z_correct<="0001110011011011";
        when 11560 => y_in <= "10101101"; x_in <= "10101000"; z_correct<="0001110010001000";
        when 11561 => y_in <= "10101101"; x_in <= "10101001"; z_correct<="0001110000110101";
        when 11562 => y_in <= "10101101"; x_in <= "10101010"; z_correct<="0001101111100010";
        when 11563 => y_in <= "10101101"; x_in <= "10101011"; z_correct<="0001101110001111";
        when 11564 => y_in <= "10101101"; x_in <= "10101100"; z_correct<="0001101100111100";
        when 11565 => y_in <= "10101101"; x_in <= "10101101"; z_correct<="0001101011101001";
        when 11566 => y_in <= "10101101"; x_in <= "10101110"; z_correct<="0001101010010110";
        when 11567 => y_in <= "10101101"; x_in <= "10101111"; z_correct<="0001101001000011";
        when 11568 => y_in <= "10101101"; x_in <= "10110000"; z_correct<="0001100111110000";
        when 11569 => y_in <= "10101101"; x_in <= "10110001"; z_correct<="0001100110011101";
        when 11570 => y_in <= "10101101"; x_in <= "10110010"; z_correct<="0001100101001010";
        when 11571 => y_in <= "10101101"; x_in <= "10110011"; z_correct<="0001100011110111";
        when 11572 => y_in <= "10101101"; x_in <= "10110100"; z_correct<="0001100010100100";
        when 11573 => y_in <= "10101101"; x_in <= "10110101"; z_correct<="0001100001010001";
        when 11574 => y_in <= "10101101"; x_in <= "10110110"; z_correct<="0001011111111110";
        when 11575 => y_in <= "10101101"; x_in <= "10110111"; z_correct<="0001011110101011";
        when 11576 => y_in <= "10101101"; x_in <= "10111000"; z_correct<="0001011101011000";
        when 11577 => y_in <= "10101101"; x_in <= "10111001"; z_correct<="0001011100000101";
        when 11578 => y_in <= "10101101"; x_in <= "10111010"; z_correct<="0001011010110010";
        when 11579 => y_in <= "10101101"; x_in <= "10111011"; z_correct<="0001011001011111";
        when 11580 => y_in <= "10101101"; x_in <= "10111100"; z_correct<="0001011000001100";
        when 11581 => y_in <= "10101101"; x_in <= "10111101"; z_correct<="0001010110111001";
        when 11582 => y_in <= "10101101"; x_in <= "10111110"; z_correct<="0001010101100110";
        when 11583 => y_in <= "10101101"; x_in <= "10111111"; z_correct<="0001010100010011";
        when 11584 => y_in <= "10101101"; x_in <= "11000000"; z_correct<="0001010011000000";
        when 11585 => y_in <= "10101101"; x_in <= "11000001"; z_correct<="0001010001101101";
        when 11586 => y_in <= "10101101"; x_in <= "11000010"; z_correct<="0001010000011010";
        when 11587 => y_in <= "10101101"; x_in <= "11000011"; z_correct<="0001001111000111";
        when 11588 => y_in <= "10101101"; x_in <= "11000100"; z_correct<="0001001101110100";
        when 11589 => y_in <= "10101101"; x_in <= "11000101"; z_correct<="0001001100100001";
        when 11590 => y_in <= "10101101"; x_in <= "11000110"; z_correct<="0001001011001110";
        when 11591 => y_in <= "10101101"; x_in <= "11000111"; z_correct<="0001001001111011";
        when 11592 => y_in <= "10101101"; x_in <= "11001000"; z_correct<="0001001000101000";
        when 11593 => y_in <= "10101101"; x_in <= "11001001"; z_correct<="0001000111010101";
        when 11594 => y_in <= "10101101"; x_in <= "11001010"; z_correct<="0001000110000010";
        when 11595 => y_in <= "10101101"; x_in <= "11001011"; z_correct<="0001000100101111";
        when 11596 => y_in <= "10101101"; x_in <= "11001100"; z_correct<="0001000011011100";
        when 11597 => y_in <= "10101101"; x_in <= "11001101"; z_correct<="0001000010001001";
        when 11598 => y_in <= "10101101"; x_in <= "11001110"; z_correct<="0001000000110110";
        when 11599 => y_in <= "10101101"; x_in <= "11001111"; z_correct<="0000111111100011";
        when 11600 => y_in <= "10101101"; x_in <= "11010000"; z_correct<="0000111110010000";
        when 11601 => y_in <= "10101101"; x_in <= "11010001"; z_correct<="0000111100111101";
        when 11602 => y_in <= "10101101"; x_in <= "11010010"; z_correct<="0000111011101010";
        when 11603 => y_in <= "10101101"; x_in <= "11010011"; z_correct<="0000111010010111";
        when 11604 => y_in <= "10101101"; x_in <= "11010100"; z_correct<="0000111001000100";
        when 11605 => y_in <= "10101101"; x_in <= "11010101"; z_correct<="0000110111110001";
        when 11606 => y_in <= "10101101"; x_in <= "11010110"; z_correct<="0000110110011110";
        when 11607 => y_in <= "10101101"; x_in <= "11010111"; z_correct<="0000110101001011";
        when 11608 => y_in <= "10101101"; x_in <= "11011000"; z_correct<="0000110011111000";
        when 11609 => y_in <= "10101101"; x_in <= "11011001"; z_correct<="0000110010100101";
        when 11610 => y_in <= "10101101"; x_in <= "11011010"; z_correct<="0000110001010010";
        when 11611 => y_in <= "10101101"; x_in <= "11011011"; z_correct<="0000101111111111";
        when 11612 => y_in <= "10101101"; x_in <= "11011100"; z_correct<="0000101110101100";
        when 11613 => y_in <= "10101101"; x_in <= "11011101"; z_correct<="0000101101011001";
        when 11614 => y_in <= "10101101"; x_in <= "11011110"; z_correct<="0000101100000110";
        when 11615 => y_in <= "10101101"; x_in <= "11011111"; z_correct<="0000101010110011";
        when 11616 => y_in <= "10101101"; x_in <= "11100000"; z_correct<="0000101001100000";
        when 11617 => y_in <= "10101101"; x_in <= "11100001"; z_correct<="0000101000001101";
        when 11618 => y_in <= "10101101"; x_in <= "11100010"; z_correct<="0000100110111010";
        when 11619 => y_in <= "10101101"; x_in <= "11100011"; z_correct<="0000100101100111";
        when 11620 => y_in <= "10101101"; x_in <= "11100100"; z_correct<="0000100100010100";
        when 11621 => y_in <= "10101101"; x_in <= "11100101"; z_correct<="0000100011000001";
        when 11622 => y_in <= "10101101"; x_in <= "11100110"; z_correct<="0000100001101110";
        when 11623 => y_in <= "10101101"; x_in <= "11100111"; z_correct<="0000100000011011";
        when 11624 => y_in <= "10101101"; x_in <= "11101000"; z_correct<="0000011111001000";
        when 11625 => y_in <= "10101101"; x_in <= "11101001"; z_correct<="0000011101110101";
        when 11626 => y_in <= "10101101"; x_in <= "11101010"; z_correct<="0000011100100010";
        when 11627 => y_in <= "10101101"; x_in <= "11101011"; z_correct<="0000011011001111";
        when 11628 => y_in <= "10101101"; x_in <= "11101100"; z_correct<="0000011001111100";
        when 11629 => y_in <= "10101101"; x_in <= "11101101"; z_correct<="0000011000101001";
        when 11630 => y_in <= "10101101"; x_in <= "11101110"; z_correct<="0000010111010110";
        when 11631 => y_in <= "10101101"; x_in <= "11101111"; z_correct<="0000010110000011";
        when 11632 => y_in <= "10101101"; x_in <= "11110000"; z_correct<="0000010100110000";
        when 11633 => y_in <= "10101101"; x_in <= "11110001"; z_correct<="0000010011011101";
        when 11634 => y_in <= "10101101"; x_in <= "11110010"; z_correct<="0000010010001010";
        when 11635 => y_in <= "10101101"; x_in <= "11110011"; z_correct<="0000010000110111";
        when 11636 => y_in <= "10101101"; x_in <= "11110100"; z_correct<="0000001111100100";
        when 11637 => y_in <= "10101101"; x_in <= "11110101"; z_correct<="0000001110010001";
        when 11638 => y_in <= "10101101"; x_in <= "11110110"; z_correct<="0000001100111110";
        when 11639 => y_in <= "10101101"; x_in <= "11110111"; z_correct<="0000001011101011";
        when 11640 => y_in <= "10101101"; x_in <= "11111000"; z_correct<="0000001010011000";
        when 11641 => y_in <= "10101101"; x_in <= "11111001"; z_correct<="0000001001000101";
        when 11642 => y_in <= "10101101"; x_in <= "11111010"; z_correct<="0000000111110010";
        when 11643 => y_in <= "10101101"; x_in <= "11111011"; z_correct<="0000000110011111";
        when 11644 => y_in <= "10101101"; x_in <= "11111100"; z_correct<="0000000101001100";
        when 11645 => y_in <= "10101101"; x_in <= "11111101"; z_correct<="0000000011111001";
        when 11646 => y_in <= "10101101"; x_in <= "11111110"; z_correct<="0000000010100110";
        when 11647 => y_in <= "10101101"; x_in <= "11111111"; z_correct<="0000000001010011";
        when 11648 => y_in <= "10101101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 11649 => y_in <= "10101101"; x_in <= "00000001"; z_correct<="1111111110101101";
        when 11650 => y_in <= "10101101"; x_in <= "00000010"; z_correct<="1111111101011010";
        when 11651 => y_in <= "10101101"; x_in <= "00000011"; z_correct<="1111111100000111";
        when 11652 => y_in <= "10101101"; x_in <= "00000100"; z_correct<="1111111010110100";
        when 11653 => y_in <= "10101101"; x_in <= "00000101"; z_correct<="1111111001100001";
        when 11654 => y_in <= "10101101"; x_in <= "00000110"; z_correct<="1111111000001110";
        when 11655 => y_in <= "10101101"; x_in <= "00000111"; z_correct<="1111110110111011";
        when 11656 => y_in <= "10101101"; x_in <= "00001000"; z_correct<="1111110101101000";
        when 11657 => y_in <= "10101101"; x_in <= "00001001"; z_correct<="1111110100010101";
        when 11658 => y_in <= "10101101"; x_in <= "00001010"; z_correct<="1111110011000010";
        when 11659 => y_in <= "10101101"; x_in <= "00001011"; z_correct<="1111110001101111";
        when 11660 => y_in <= "10101101"; x_in <= "00001100"; z_correct<="1111110000011100";
        when 11661 => y_in <= "10101101"; x_in <= "00001101"; z_correct<="1111101111001001";
        when 11662 => y_in <= "10101101"; x_in <= "00001110"; z_correct<="1111101101110110";
        when 11663 => y_in <= "10101101"; x_in <= "00001111"; z_correct<="1111101100100011";
        when 11664 => y_in <= "10101101"; x_in <= "00010000"; z_correct<="1111101011010000";
        when 11665 => y_in <= "10101101"; x_in <= "00010001"; z_correct<="1111101001111101";
        when 11666 => y_in <= "10101101"; x_in <= "00010010"; z_correct<="1111101000101010";
        when 11667 => y_in <= "10101101"; x_in <= "00010011"; z_correct<="1111100111010111";
        when 11668 => y_in <= "10101101"; x_in <= "00010100"; z_correct<="1111100110000100";
        when 11669 => y_in <= "10101101"; x_in <= "00010101"; z_correct<="1111100100110001";
        when 11670 => y_in <= "10101101"; x_in <= "00010110"; z_correct<="1111100011011110";
        when 11671 => y_in <= "10101101"; x_in <= "00010111"; z_correct<="1111100010001011";
        when 11672 => y_in <= "10101101"; x_in <= "00011000"; z_correct<="1111100000111000";
        when 11673 => y_in <= "10101101"; x_in <= "00011001"; z_correct<="1111011111100101";
        when 11674 => y_in <= "10101101"; x_in <= "00011010"; z_correct<="1111011110010010";
        when 11675 => y_in <= "10101101"; x_in <= "00011011"; z_correct<="1111011100111111";
        when 11676 => y_in <= "10101101"; x_in <= "00011100"; z_correct<="1111011011101100";
        when 11677 => y_in <= "10101101"; x_in <= "00011101"; z_correct<="1111011010011001";
        when 11678 => y_in <= "10101101"; x_in <= "00011110"; z_correct<="1111011001000110";
        when 11679 => y_in <= "10101101"; x_in <= "00011111"; z_correct<="1111010111110011";
        when 11680 => y_in <= "10101101"; x_in <= "00100000"; z_correct<="1111010110100000";
        when 11681 => y_in <= "10101101"; x_in <= "00100001"; z_correct<="1111010101001101";
        when 11682 => y_in <= "10101101"; x_in <= "00100010"; z_correct<="1111010011111010";
        when 11683 => y_in <= "10101101"; x_in <= "00100011"; z_correct<="1111010010100111";
        when 11684 => y_in <= "10101101"; x_in <= "00100100"; z_correct<="1111010001010100";
        when 11685 => y_in <= "10101101"; x_in <= "00100101"; z_correct<="1111010000000001";
        when 11686 => y_in <= "10101101"; x_in <= "00100110"; z_correct<="1111001110101110";
        when 11687 => y_in <= "10101101"; x_in <= "00100111"; z_correct<="1111001101011011";
        when 11688 => y_in <= "10101101"; x_in <= "00101000"; z_correct<="1111001100001000";
        when 11689 => y_in <= "10101101"; x_in <= "00101001"; z_correct<="1111001010110101";
        when 11690 => y_in <= "10101101"; x_in <= "00101010"; z_correct<="1111001001100010";
        when 11691 => y_in <= "10101101"; x_in <= "00101011"; z_correct<="1111001000001111";
        when 11692 => y_in <= "10101101"; x_in <= "00101100"; z_correct<="1111000110111100";
        when 11693 => y_in <= "10101101"; x_in <= "00101101"; z_correct<="1111000101101001";
        when 11694 => y_in <= "10101101"; x_in <= "00101110"; z_correct<="1111000100010110";
        when 11695 => y_in <= "10101101"; x_in <= "00101111"; z_correct<="1111000011000011";
        when 11696 => y_in <= "10101101"; x_in <= "00110000"; z_correct<="1111000001110000";
        when 11697 => y_in <= "10101101"; x_in <= "00110001"; z_correct<="1111000000011101";
        when 11698 => y_in <= "10101101"; x_in <= "00110010"; z_correct<="1110111111001010";
        when 11699 => y_in <= "10101101"; x_in <= "00110011"; z_correct<="1110111101110111";
        when 11700 => y_in <= "10101101"; x_in <= "00110100"; z_correct<="1110111100100100";
        when 11701 => y_in <= "10101101"; x_in <= "00110101"; z_correct<="1110111011010001";
        when 11702 => y_in <= "10101101"; x_in <= "00110110"; z_correct<="1110111001111110";
        when 11703 => y_in <= "10101101"; x_in <= "00110111"; z_correct<="1110111000101011";
        when 11704 => y_in <= "10101101"; x_in <= "00111000"; z_correct<="1110110111011000";
        when 11705 => y_in <= "10101101"; x_in <= "00111001"; z_correct<="1110110110000101";
        when 11706 => y_in <= "10101101"; x_in <= "00111010"; z_correct<="1110110100110010";
        when 11707 => y_in <= "10101101"; x_in <= "00111011"; z_correct<="1110110011011111";
        when 11708 => y_in <= "10101101"; x_in <= "00111100"; z_correct<="1110110010001100";
        when 11709 => y_in <= "10101101"; x_in <= "00111101"; z_correct<="1110110000111001";
        when 11710 => y_in <= "10101101"; x_in <= "00111110"; z_correct<="1110101111100110";
        when 11711 => y_in <= "10101101"; x_in <= "00111111"; z_correct<="1110101110010011";
        when 11712 => y_in <= "10101101"; x_in <= "01000000"; z_correct<="1110101101000000";
        when 11713 => y_in <= "10101101"; x_in <= "01000001"; z_correct<="1110101011101101";
        when 11714 => y_in <= "10101101"; x_in <= "01000010"; z_correct<="1110101010011010";
        when 11715 => y_in <= "10101101"; x_in <= "01000011"; z_correct<="1110101001000111";
        when 11716 => y_in <= "10101101"; x_in <= "01000100"; z_correct<="1110100111110100";
        when 11717 => y_in <= "10101101"; x_in <= "01000101"; z_correct<="1110100110100001";
        when 11718 => y_in <= "10101101"; x_in <= "01000110"; z_correct<="1110100101001110";
        when 11719 => y_in <= "10101101"; x_in <= "01000111"; z_correct<="1110100011111011";
        when 11720 => y_in <= "10101101"; x_in <= "01001000"; z_correct<="1110100010101000";
        when 11721 => y_in <= "10101101"; x_in <= "01001001"; z_correct<="1110100001010101";
        when 11722 => y_in <= "10101101"; x_in <= "01001010"; z_correct<="1110100000000010";
        when 11723 => y_in <= "10101101"; x_in <= "01001011"; z_correct<="1110011110101111";
        when 11724 => y_in <= "10101101"; x_in <= "01001100"; z_correct<="1110011101011100";
        when 11725 => y_in <= "10101101"; x_in <= "01001101"; z_correct<="1110011100001001";
        when 11726 => y_in <= "10101101"; x_in <= "01001110"; z_correct<="1110011010110110";
        when 11727 => y_in <= "10101101"; x_in <= "01001111"; z_correct<="1110011001100011";
        when 11728 => y_in <= "10101101"; x_in <= "01010000"; z_correct<="1110011000010000";
        when 11729 => y_in <= "10101101"; x_in <= "01010001"; z_correct<="1110010110111101";
        when 11730 => y_in <= "10101101"; x_in <= "01010010"; z_correct<="1110010101101010";
        when 11731 => y_in <= "10101101"; x_in <= "01010011"; z_correct<="1110010100010111";
        when 11732 => y_in <= "10101101"; x_in <= "01010100"; z_correct<="1110010011000100";
        when 11733 => y_in <= "10101101"; x_in <= "01010101"; z_correct<="1110010001110001";
        when 11734 => y_in <= "10101101"; x_in <= "01010110"; z_correct<="1110010000011110";
        when 11735 => y_in <= "10101101"; x_in <= "01010111"; z_correct<="1110001111001011";
        when 11736 => y_in <= "10101101"; x_in <= "01011000"; z_correct<="1110001101111000";
        when 11737 => y_in <= "10101101"; x_in <= "01011001"; z_correct<="1110001100100101";
        when 11738 => y_in <= "10101101"; x_in <= "01011010"; z_correct<="1110001011010010";
        when 11739 => y_in <= "10101101"; x_in <= "01011011"; z_correct<="1110001001111111";
        when 11740 => y_in <= "10101101"; x_in <= "01011100"; z_correct<="1110001000101100";
        when 11741 => y_in <= "10101101"; x_in <= "01011101"; z_correct<="1110000111011001";
        when 11742 => y_in <= "10101101"; x_in <= "01011110"; z_correct<="1110000110000110";
        when 11743 => y_in <= "10101101"; x_in <= "01011111"; z_correct<="1110000100110011";
        when 11744 => y_in <= "10101101"; x_in <= "01100000"; z_correct<="1110000011100000";
        when 11745 => y_in <= "10101101"; x_in <= "01100001"; z_correct<="1110000010001101";
        when 11746 => y_in <= "10101101"; x_in <= "01100010"; z_correct<="1110000000111010";
        when 11747 => y_in <= "10101101"; x_in <= "01100011"; z_correct<="1101111111100111";
        when 11748 => y_in <= "10101101"; x_in <= "01100100"; z_correct<="1101111110010100";
        when 11749 => y_in <= "10101101"; x_in <= "01100101"; z_correct<="1101111101000001";
        when 11750 => y_in <= "10101101"; x_in <= "01100110"; z_correct<="1101111011101110";
        when 11751 => y_in <= "10101101"; x_in <= "01100111"; z_correct<="1101111010011011";
        when 11752 => y_in <= "10101101"; x_in <= "01101000"; z_correct<="1101111001001000";
        when 11753 => y_in <= "10101101"; x_in <= "01101001"; z_correct<="1101110111110101";
        when 11754 => y_in <= "10101101"; x_in <= "01101010"; z_correct<="1101110110100010";
        when 11755 => y_in <= "10101101"; x_in <= "01101011"; z_correct<="1101110101001111";
        when 11756 => y_in <= "10101101"; x_in <= "01101100"; z_correct<="1101110011111100";
        when 11757 => y_in <= "10101101"; x_in <= "01101101"; z_correct<="1101110010101001";
        when 11758 => y_in <= "10101101"; x_in <= "01101110"; z_correct<="1101110001010110";
        when 11759 => y_in <= "10101101"; x_in <= "01101111"; z_correct<="1101110000000011";
        when 11760 => y_in <= "10101101"; x_in <= "01110000"; z_correct<="1101101110110000";
        when 11761 => y_in <= "10101101"; x_in <= "01110001"; z_correct<="1101101101011101";
        when 11762 => y_in <= "10101101"; x_in <= "01110010"; z_correct<="1101101100001010";
        when 11763 => y_in <= "10101101"; x_in <= "01110011"; z_correct<="1101101010110111";
        when 11764 => y_in <= "10101101"; x_in <= "01110100"; z_correct<="1101101001100100";
        when 11765 => y_in <= "10101101"; x_in <= "01110101"; z_correct<="1101101000010001";
        when 11766 => y_in <= "10101101"; x_in <= "01110110"; z_correct<="1101100110111110";
        when 11767 => y_in <= "10101101"; x_in <= "01110111"; z_correct<="1101100101101011";
        when 11768 => y_in <= "10101101"; x_in <= "01111000"; z_correct<="1101100100011000";
        when 11769 => y_in <= "10101101"; x_in <= "01111001"; z_correct<="1101100011000101";
        when 11770 => y_in <= "10101101"; x_in <= "01111010"; z_correct<="1101100001110010";
        when 11771 => y_in <= "10101101"; x_in <= "01111011"; z_correct<="1101100000011111";
        when 11772 => y_in <= "10101101"; x_in <= "01111100"; z_correct<="1101011111001100";
        when 11773 => y_in <= "10101101"; x_in <= "01111101"; z_correct<="1101011101111001";
        when 11774 => y_in <= "10101101"; x_in <= "01111110"; z_correct<="1101011100100110";
        when 11775 => y_in <= "10101101"; x_in <= "01111111"; z_correct<="1101011011010011";
        when 11776 => y_in <= "10101110"; x_in <= "10000000"; z_correct<="0010100100000000";
        when 11777 => y_in <= "10101110"; x_in <= "10000001"; z_correct<="0010100010101110";
        when 11778 => y_in <= "10101110"; x_in <= "10000010"; z_correct<="0010100001011100";
        when 11779 => y_in <= "10101110"; x_in <= "10000011"; z_correct<="0010100000001010";
        when 11780 => y_in <= "10101110"; x_in <= "10000100"; z_correct<="0010011110111000";
        when 11781 => y_in <= "10101110"; x_in <= "10000101"; z_correct<="0010011101100110";
        when 11782 => y_in <= "10101110"; x_in <= "10000110"; z_correct<="0010011100010100";
        when 11783 => y_in <= "10101110"; x_in <= "10000111"; z_correct<="0010011011000010";
        when 11784 => y_in <= "10101110"; x_in <= "10001000"; z_correct<="0010011001110000";
        when 11785 => y_in <= "10101110"; x_in <= "10001001"; z_correct<="0010011000011110";
        when 11786 => y_in <= "10101110"; x_in <= "10001010"; z_correct<="0010010111001100";
        when 11787 => y_in <= "10101110"; x_in <= "10001011"; z_correct<="0010010101111010";
        when 11788 => y_in <= "10101110"; x_in <= "10001100"; z_correct<="0010010100101000";
        when 11789 => y_in <= "10101110"; x_in <= "10001101"; z_correct<="0010010011010110";
        when 11790 => y_in <= "10101110"; x_in <= "10001110"; z_correct<="0010010010000100";
        when 11791 => y_in <= "10101110"; x_in <= "10001111"; z_correct<="0010010000110010";
        when 11792 => y_in <= "10101110"; x_in <= "10010000"; z_correct<="0010001111100000";
        when 11793 => y_in <= "10101110"; x_in <= "10010001"; z_correct<="0010001110001110";
        when 11794 => y_in <= "10101110"; x_in <= "10010010"; z_correct<="0010001100111100";
        when 11795 => y_in <= "10101110"; x_in <= "10010011"; z_correct<="0010001011101010";
        when 11796 => y_in <= "10101110"; x_in <= "10010100"; z_correct<="0010001010011000";
        when 11797 => y_in <= "10101110"; x_in <= "10010101"; z_correct<="0010001001000110";
        when 11798 => y_in <= "10101110"; x_in <= "10010110"; z_correct<="0010000111110100";
        when 11799 => y_in <= "10101110"; x_in <= "10010111"; z_correct<="0010000110100010";
        when 11800 => y_in <= "10101110"; x_in <= "10011000"; z_correct<="0010000101010000";
        when 11801 => y_in <= "10101110"; x_in <= "10011001"; z_correct<="0010000011111110";
        when 11802 => y_in <= "10101110"; x_in <= "10011010"; z_correct<="0010000010101100";
        when 11803 => y_in <= "10101110"; x_in <= "10011011"; z_correct<="0010000001011010";
        when 11804 => y_in <= "10101110"; x_in <= "10011100"; z_correct<="0010000000001000";
        when 11805 => y_in <= "10101110"; x_in <= "10011101"; z_correct<="0001111110110110";
        when 11806 => y_in <= "10101110"; x_in <= "10011110"; z_correct<="0001111101100100";
        when 11807 => y_in <= "10101110"; x_in <= "10011111"; z_correct<="0001111100010010";
        when 11808 => y_in <= "10101110"; x_in <= "10100000"; z_correct<="0001111011000000";
        when 11809 => y_in <= "10101110"; x_in <= "10100001"; z_correct<="0001111001101110";
        when 11810 => y_in <= "10101110"; x_in <= "10100010"; z_correct<="0001111000011100";
        when 11811 => y_in <= "10101110"; x_in <= "10100011"; z_correct<="0001110111001010";
        when 11812 => y_in <= "10101110"; x_in <= "10100100"; z_correct<="0001110101111000";
        when 11813 => y_in <= "10101110"; x_in <= "10100101"; z_correct<="0001110100100110";
        when 11814 => y_in <= "10101110"; x_in <= "10100110"; z_correct<="0001110011010100";
        when 11815 => y_in <= "10101110"; x_in <= "10100111"; z_correct<="0001110010000010";
        when 11816 => y_in <= "10101110"; x_in <= "10101000"; z_correct<="0001110000110000";
        when 11817 => y_in <= "10101110"; x_in <= "10101001"; z_correct<="0001101111011110";
        when 11818 => y_in <= "10101110"; x_in <= "10101010"; z_correct<="0001101110001100";
        when 11819 => y_in <= "10101110"; x_in <= "10101011"; z_correct<="0001101100111010";
        when 11820 => y_in <= "10101110"; x_in <= "10101100"; z_correct<="0001101011101000";
        when 11821 => y_in <= "10101110"; x_in <= "10101101"; z_correct<="0001101010010110";
        when 11822 => y_in <= "10101110"; x_in <= "10101110"; z_correct<="0001101001000100";
        when 11823 => y_in <= "10101110"; x_in <= "10101111"; z_correct<="0001100111110010";
        when 11824 => y_in <= "10101110"; x_in <= "10110000"; z_correct<="0001100110100000";
        when 11825 => y_in <= "10101110"; x_in <= "10110001"; z_correct<="0001100101001110";
        when 11826 => y_in <= "10101110"; x_in <= "10110010"; z_correct<="0001100011111100";
        when 11827 => y_in <= "10101110"; x_in <= "10110011"; z_correct<="0001100010101010";
        when 11828 => y_in <= "10101110"; x_in <= "10110100"; z_correct<="0001100001011000";
        when 11829 => y_in <= "10101110"; x_in <= "10110101"; z_correct<="0001100000000110";
        when 11830 => y_in <= "10101110"; x_in <= "10110110"; z_correct<="0001011110110100";
        when 11831 => y_in <= "10101110"; x_in <= "10110111"; z_correct<="0001011101100010";
        when 11832 => y_in <= "10101110"; x_in <= "10111000"; z_correct<="0001011100010000";
        when 11833 => y_in <= "10101110"; x_in <= "10111001"; z_correct<="0001011010111110";
        when 11834 => y_in <= "10101110"; x_in <= "10111010"; z_correct<="0001011001101100";
        when 11835 => y_in <= "10101110"; x_in <= "10111011"; z_correct<="0001011000011010";
        when 11836 => y_in <= "10101110"; x_in <= "10111100"; z_correct<="0001010111001000";
        when 11837 => y_in <= "10101110"; x_in <= "10111101"; z_correct<="0001010101110110";
        when 11838 => y_in <= "10101110"; x_in <= "10111110"; z_correct<="0001010100100100";
        when 11839 => y_in <= "10101110"; x_in <= "10111111"; z_correct<="0001010011010010";
        when 11840 => y_in <= "10101110"; x_in <= "11000000"; z_correct<="0001010010000000";
        when 11841 => y_in <= "10101110"; x_in <= "11000001"; z_correct<="0001010000101110";
        when 11842 => y_in <= "10101110"; x_in <= "11000010"; z_correct<="0001001111011100";
        when 11843 => y_in <= "10101110"; x_in <= "11000011"; z_correct<="0001001110001010";
        when 11844 => y_in <= "10101110"; x_in <= "11000100"; z_correct<="0001001100111000";
        when 11845 => y_in <= "10101110"; x_in <= "11000101"; z_correct<="0001001011100110";
        when 11846 => y_in <= "10101110"; x_in <= "11000110"; z_correct<="0001001010010100";
        when 11847 => y_in <= "10101110"; x_in <= "11000111"; z_correct<="0001001001000010";
        when 11848 => y_in <= "10101110"; x_in <= "11001000"; z_correct<="0001000111110000";
        when 11849 => y_in <= "10101110"; x_in <= "11001001"; z_correct<="0001000110011110";
        when 11850 => y_in <= "10101110"; x_in <= "11001010"; z_correct<="0001000101001100";
        when 11851 => y_in <= "10101110"; x_in <= "11001011"; z_correct<="0001000011111010";
        when 11852 => y_in <= "10101110"; x_in <= "11001100"; z_correct<="0001000010101000";
        when 11853 => y_in <= "10101110"; x_in <= "11001101"; z_correct<="0001000001010110";
        when 11854 => y_in <= "10101110"; x_in <= "11001110"; z_correct<="0001000000000100";
        when 11855 => y_in <= "10101110"; x_in <= "11001111"; z_correct<="0000111110110010";
        when 11856 => y_in <= "10101110"; x_in <= "11010000"; z_correct<="0000111101100000";
        when 11857 => y_in <= "10101110"; x_in <= "11010001"; z_correct<="0000111100001110";
        when 11858 => y_in <= "10101110"; x_in <= "11010010"; z_correct<="0000111010111100";
        when 11859 => y_in <= "10101110"; x_in <= "11010011"; z_correct<="0000111001101010";
        when 11860 => y_in <= "10101110"; x_in <= "11010100"; z_correct<="0000111000011000";
        when 11861 => y_in <= "10101110"; x_in <= "11010101"; z_correct<="0000110111000110";
        when 11862 => y_in <= "10101110"; x_in <= "11010110"; z_correct<="0000110101110100";
        when 11863 => y_in <= "10101110"; x_in <= "11010111"; z_correct<="0000110100100010";
        when 11864 => y_in <= "10101110"; x_in <= "11011000"; z_correct<="0000110011010000";
        when 11865 => y_in <= "10101110"; x_in <= "11011001"; z_correct<="0000110001111110";
        when 11866 => y_in <= "10101110"; x_in <= "11011010"; z_correct<="0000110000101100";
        when 11867 => y_in <= "10101110"; x_in <= "11011011"; z_correct<="0000101111011010";
        when 11868 => y_in <= "10101110"; x_in <= "11011100"; z_correct<="0000101110001000";
        when 11869 => y_in <= "10101110"; x_in <= "11011101"; z_correct<="0000101100110110";
        when 11870 => y_in <= "10101110"; x_in <= "11011110"; z_correct<="0000101011100100";
        when 11871 => y_in <= "10101110"; x_in <= "11011111"; z_correct<="0000101010010010";
        when 11872 => y_in <= "10101110"; x_in <= "11100000"; z_correct<="0000101001000000";
        when 11873 => y_in <= "10101110"; x_in <= "11100001"; z_correct<="0000100111101110";
        when 11874 => y_in <= "10101110"; x_in <= "11100010"; z_correct<="0000100110011100";
        when 11875 => y_in <= "10101110"; x_in <= "11100011"; z_correct<="0000100101001010";
        when 11876 => y_in <= "10101110"; x_in <= "11100100"; z_correct<="0000100011111000";
        when 11877 => y_in <= "10101110"; x_in <= "11100101"; z_correct<="0000100010100110";
        when 11878 => y_in <= "10101110"; x_in <= "11100110"; z_correct<="0000100001010100";
        when 11879 => y_in <= "10101110"; x_in <= "11100111"; z_correct<="0000100000000010";
        when 11880 => y_in <= "10101110"; x_in <= "11101000"; z_correct<="0000011110110000";
        when 11881 => y_in <= "10101110"; x_in <= "11101001"; z_correct<="0000011101011110";
        when 11882 => y_in <= "10101110"; x_in <= "11101010"; z_correct<="0000011100001100";
        when 11883 => y_in <= "10101110"; x_in <= "11101011"; z_correct<="0000011010111010";
        when 11884 => y_in <= "10101110"; x_in <= "11101100"; z_correct<="0000011001101000";
        when 11885 => y_in <= "10101110"; x_in <= "11101101"; z_correct<="0000011000010110";
        when 11886 => y_in <= "10101110"; x_in <= "11101110"; z_correct<="0000010111000100";
        when 11887 => y_in <= "10101110"; x_in <= "11101111"; z_correct<="0000010101110010";
        when 11888 => y_in <= "10101110"; x_in <= "11110000"; z_correct<="0000010100100000";
        when 11889 => y_in <= "10101110"; x_in <= "11110001"; z_correct<="0000010011001110";
        when 11890 => y_in <= "10101110"; x_in <= "11110010"; z_correct<="0000010001111100";
        when 11891 => y_in <= "10101110"; x_in <= "11110011"; z_correct<="0000010000101010";
        when 11892 => y_in <= "10101110"; x_in <= "11110100"; z_correct<="0000001111011000";
        when 11893 => y_in <= "10101110"; x_in <= "11110101"; z_correct<="0000001110000110";
        when 11894 => y_in <= "10101110"; x_in <= "11110110"; z_correct<="0000001100110100";
        when 11895 => y_in <= "10101110"; x_in <= "11110111"; z_correct<="0000001011100010";
        when 11896 => y_in <= "10101110"; x_in <= "11111000"; z_correct<="0000001010010000";
        when 11897 => y_in <= "10101110"; x_in <= "11111001"; z_correct<="0000001000111110";
        when 11898 => y_in <= "10101110"; x_in <= "11111010"; z_correct<="0000000111101100";
        when 11899 => y_in <= "10101110"; x_in <= "11111011"; z_correct<="0000000110011010";
        when 11900 => y_in <= "10101110"; x_in <= "11111100"; z_correct<="0000000101001000";
        when 11901 => y_in <= "10101110"; x_in <= "11111101"; z_correct<="0000000011110110";
        when 11902 => y_in <= "10101110"; x_in <= "11111110"; z_correct<="0000000010100100";
        when 11903 => y_in <= "10101110"; x_in <= "11111111"; z_correct<="0000000001010010";
        when 11904 => y_in <= "10101110"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 11905 => y_in <= "10101110"; x_in <= "00000001"; z_correct<="1111111110101110";
        when 11906 => y_in <= "10101110"; x_in <= "00000010"; z_correct<="1111111101011100";
        when 11907 => y_in <= "10101110"; x_in <= "00000011"; z_correct<="1111111100001010";
        when 11908 => y_in <= "10101110"; x_in <= "00000100"; z_correct<="1111111010111000";
        when 11909 => y_in <= "10101110"; x_in <= "00000101"; z_correct<="1111111001100110";
        when 11910 => y_in <= "10101110"; x_in <= "00000110"; z_correct<="1111111000010100";
        when 11911 => y_in <= "10101110"; x_in <= "00000111"; z_correct<="1111110111000010";
        when 11912 => y_in <= "10101110"; x_in <= "00001000"; z_correct<="1111110101110000";
        when 11913 => y_in <= "10101110"; x_in <= "00001001"; z_correct<="1111110100011110";
        when 11914 => y_in <= "10101110"; x_in <= "00001010"; z_correct<="1111110011001100";
        when 11915 => y_in <= "10101110"; x_in <= "00001011"; z_correct<="1111110001111010";
        when 11916 => y_in <= "10101110"; x_in <= "00001100"; z_correct<="1111110000101000";
        when 11917 => y_in <= "10101110"; x_in <= "00001101"; z_correct<="1111101111010110";
        when 11918 => y_in <= "10101110"; x_in <= "00001110"; z_correct<="1111101110000100";
        when 11919 => y_in <= "10101110"; x_in <= "00001111"; z_correct<="1111101100110010";
        when 11920 => y_in <= "10101110"; x_in <= "00010000"; z_correct<="1111101011100000";
        when 11921 => y_in <= "10101110"; x_in <= "00010001"; z_correct<="1111101010001110";
        when 11922 => y_in <= "10101110"; x_in <= "00010010"; z_correct<="1111101000111100";
        when 11923 => y_in <= "10101110"; x_in <= "00010011"; z_correct<="1111100111101010";
        when 11924 => y_in <= "10101110"; x_in <= "00010100"; z_correct<="1111100110011000";
        when 11925 => y_in <= "10101110"; x_in <= "00010101"; z_correct<="1111100101000110";
        when 11926 => y_in <= "10101110"; x_in <= "00010110"; z_correct<="1111100011110100";
        when 11927 => y_in <= "10101110"; x_in <= "00010111"; z_correct<="1111100010100010";
        when 11928 => y_in <= "10101110"; x_in <= "00011000"; z_correct<="1111100001010000";
        when 11929 => y_in <= "10101110"; x_in <= "00011001"; z_correct<="1111011111111110";
        when 11930 => y_in <= "10101110"; x_in <= "00011010"; z_correct<="1111011110101100";
        when 11931 => y_in <= "10101110"; x_in <= "00011011"; z_correct<="1111011101011010";
        when 11932 => y_in <= "10101110"; x_in <= "00011100"; z_correct<="1111011100001000";
        when 11933 => y_in <= "10101110"; x_in <= "00011101"; z_correct<="1111011010110110";
        when 11934 => y_in <= "10101110"; x_in <= "00011110"; z_correct<="1111011001100100";
        when 11935 => y_in <= "10101110"; x_in <= "00011111"; z_correct<="1111011000010010";
        when 11936 => y_in <= "10101110"; x_in <= "00100000"; z_correct<="1111010111000000";
        when 11937 => y_in <= "10101110"; x_in <= "00100001"; z_correct<="1111010101101110";
        when 11938 => y_in <= "10101110"; x_in <= "00100010"; z_correct<="1111010100011100";
        when 11939 => y_in <= "10101110"; x_in <= "00100011"; z_correct<="1111010011001010";
        when 11940 => y_in <= "10101110"; x_in <= "00100100"; z_correct<="1111010001111000";
        when 11941 => y_in <= "10101110"; x_in <= "00100101"; z_correct<="1111010000100110";
        when 11942 => y_in <= "10101110"; x_in <= "00100110"; z_correct<="1111001111010100";
        when 11943 => y_in <= "10101110"; x_in <= "00100111"; z_correct<="1111001110000010";
        when 11944 => y_in <= "10101110"; x_in <= "00101000"; z_correct<="1111001100110000";
        when 11945 => y_in <= "10101110"; x_in <= "00101001"; z_correct<="1111001011011110";
        when 11946 => y_in <= "10101110"; x_in <= "00101010"; z_correct<="1111001010001100";
        when 11947 => y_in <= "10101110"; x_in <= "00101011"; z_correct<="1111001000111010";
        when 11948 => y_in <= "10101110"; x_in <= "00101100"; z_correct<="1111000111101000";
        when 11949 => y_in <= "10101110"; x_in <= "00101101"; z_correct<="1111000110010110";
        when 11950 => y_in <= "10101110"; x_in <= "00101110"; z_correct<="1111000101000100";
        when 11951 => y_in <= "10101110"; x_in <= "00101111"; z_correct<="1111000011110010";
        when 11952 => y_in <= "10101110"; x_in <= "00110000"; z_correct<="1111000010100000";
        when 11953 => y_in <= "10101110"; x_in <= "00110001"; z_correct<="1111000001001110";
        when 11954 => y_in <= "10101110"; x_in <= "00110010"; z_correct<="1110111111111100";
        when 11955 => y_in <= "10101110"; x_in <= "00110011"; z_correct<="1110111110101010";
        when 11956 => y_in <= "10101110"; x_in <= "00110100"; z_correct<="1110111101011000";
        when 11957 => y_in <= "10101110"; x_in <= "00110101"; z_correct<="1110111100000110";
        when 11958 => y_in <= "10101110"; x_in <= "00110110"; z_correct<="1110111010110100";
        when 11959 => y_in <= "10101110"; x_in <= "00110111"; z_correct<="1110111001100010";
        when 11960 => y_in <= "10101110"; x_in <= "00111000"; z_correct<="1110111000010000";
        when 11961 => y_in <= "10101110"; x_in <= "00111001"; z_correct<="1110110110111110";
        when 11962 => y_in <= "10101110"; x_in <= "00111010"; z_correct<="1110110101101100";
        when 11963 => y_in <= "10101110"; x_in <= "00111011"; z_correct<="1110110100011010";
        when 11964 => y_in <= "10101110"; x_in <= "00111100"; z_correct<="1110110011001000";
        when 11965 => y_in <= "10101110"; x_in <= "00111101"; z_correct<="1110110001110110";
        when 11966 => y_in <= "10101110"; x_in <= "00111110"; z_correct<="1110110000100100";
        when 11967 => y_in <= "10101110"; x_in <= "00111111"; z_correct<="1110101111010010";
        when 11968 => y_in <= "10101110"; x_in <= "01000000"; z_correct<="1110101110000000";
        when 11969 => y_in <= "10101110"; x_in <= "01000001"; z_correct<="1110101100101110";
        when 11970 => y_in <= "10101110"; x_in <= "01000010"; z_correct<="1110101011011100";
        when 11971 => y_in <= "10101110"; x_in <= "01000011"; z_correct<="1110101010001010";
        when 11972 => y_in <= "10101110"; x_in <= "01000100"; z_correct<="1110101000111000";
        when 11973 => y_in <= "10101110"; x_in <= "01000101"; z_correct<="1110100111100110";
        when 11974 => y_in <= "10101110"; x_in <= "01000110"; z_correct<="1110100110010100";
        when 11975 => y_in <= "10101110"; x_in <= "01000111"; z_correct<="1110100101000010";
        when 11976 => y_in <= "10101110"; x_in <= "01001000"; z_correct<="1110100011110000";
        when 11977 => y_in <= "10101110"; x_in <= "01001001"; z_correct<="1110100010011110";
        when 11978 => y_in <= "10101110"; x_in <= "01001010"; z_correct<="1110100001001100";
        when 11979 => y_in <= "10101110"; x_in <= "01001011"; z_correct<="1110011111111010";
        when 11980 => y_in <= "10101110"; x_in <= "01001100"; z_correct<="1110011110101000";
        when 11981 => y_in <= "10101110"; x_in <= "01001101"; z_correct<="1110011101010110";
        when 11982 => y_in <= "10101110"; x_in <= "01001110"; z_correct<="1110011100000100";
        when 11983 => y_in <= "10101110"; x_in <= "01001111"; z_correct<="1110011010110010";
        when 11984 => y_in <= "10101110"; x_in <= "01010000"; z_correct<="1110011001100000";
        when 11985 => y_in <= "10101110"; x_in <= "01010001"; z_correct<="1110011000001110";
        when 11986 => y_in <= "10101110"; x_in <= "01010010"; z_correct<="1110010110111100";
        when 11987 => y_in <= "10101110"; x_in <= "01010011"; z_correct<="1110010101101010";
        when 11988 => y_in <= "10101110"; x_in <= "01010100"; z_correct<="1110010100011000";
        when 11989 => y_in <= "10101110"; x_in <= "01010101"; z_correct<="1110010011000110";
        when 11990 => y_in <= "10101110"; x_in <= "01010110"; z_correct<="1110010001110100";
        when 11991 => y_in <= "10101110"; x_in <= "01010111"; z_correct<="1110010000100010";
        when 11992 => y_in <= "10101110"; x_in <= "01011000"; z_correct<="1110001111010000";
        when 11993 => y_in <= "10101110"; x_in <= "01011001"; z_correct<="1110001101111110";
        when 11994 => y_in <= "10101110"; x_in <= "01011010"; z_correct<="1110001100101100";
        when 11995 => y_in <= "10101110"; x_in <= "01011011"; z_correct<="1110001011011010";
        when 11996 => y_in <= "10101110"; x_in <= "01011100"; z_correct<="1110001010001000";
        when 11997 => y_in <= "10101110"; x_in <= "01011101"; z_correct<="1110001000110110";
        when 11998 => y_in <= "10101110"; x_in <= "01011110"; z_correct<="1110000111100100";
        when 11999 => y_in <= "10101110"; x_in <= "01011111"; z_correct<="1110000110010010";
        when 12000 => y_in <= "10101110"; x_in <= "01100000"; z_correct<="1110000101000000";
        when 12001 => y_in <= "10101110"; x_in <= "01100001"; z_correct<="1110000011101110";
        when 12002 => y_in <= "10101110"; x_in <= "01100010"; z_correct<="1110000010011100";
        when 12003 => y_in <= "10101110"; x_in <= "01100011"; z_correct<="1110000001001010";
        when 12004 => y_in <= "10101110"; x_in <= "01100100"; z_correct<="1101111111111000";
        when 12005 => y_in <= "10101110"; x_in <= "01100101"; z_correct<="1101111110100110";
        when 12006 => y_in <= "10101110"; x_in <= "01100110"; z_correct<="1101111101010100";
        when 12007 => y_in <= "10101110"; x_in <= "01100111"; z_correct<="1101111100000010";
        when 12008 => y_in <= "10101110"; x_in <= "01101000"; z_correct<="1101111010110000";
        when 12009 => y_in <= "10101110"; x_in <= "01101001"; z_correct<="1101111001011110";
        when 12010 => y_in <= "10101110"; x_in <= "01101010"; z_correct<="1101111000001100";
        when 12011 => y_in <= "10101110"; x_in <= "01101011"; z_correct<="1101110110111010";
        when 12012 => y_in <= "10101110"; x_in <= "01101100"; z_correct<="1101110101101000";
        when 12013 => y_in <= "10101110"; x_in <= "01101101"; z_correct<="1101110100010110";
        when 12014 => y_in <= "10101110"; x_in <= "01101110"; z_correct<="1101110011000100";
        when 12015 => y_in <= "10101110"; x_in <= "01101111"; z_correct<="1101110001110010";
        when 12016 => y_in <= "10101110"; x_in <= "01110000"; z_correct<="1101110000100000";
        when 12017 => y_in <= "10101110"; x_in <= "01110001"; z_correct<="1101101111001110";
        when 12018 => y_in <= "10101110"; x_in <= "01110010"; z_correct<="1101101101111100";
        when 12019 => y_in <= "10101110"; x_in <= "01110011"; z_correct<="1101101100101010";
        when 12020 => y_in <= "10101110"; x_in <= "01110100"; z_correct<="1101101011011000";
        when 12021 => y_in <= "10101110"; x_in <= "01110101"; z_correct<="1101101010000110";
        when 12022 => y_in <= "10101110"; x_in <= "01110110"; z_correct<="1101101000110100";
        when 12023 => y_in <= "10101110"; x_in <= "01110111"; z_correct<="1101100111100010";
        when 12024 => y_in <= "10101110"; x_in <= "01111000"; z_correct<="1101100110010000";
        when 12025 => y_in <= "10101110"; x_in <= "01111001"; z_correct<="1101100100111110";
        when 12026 => y_in <= "10101110"; x_in <= "01111010"; z_correct<="1101100011101100";
        when 12027 => y_in <= "10101110"; x_in <= "01111011"; z_correct<="1101100010011010";
        when 12028 => y_in <= "10101110"; x_in <= "01111100"; z_correct<="1101100001001000";
        when 12029 => y_in <= "10101110"; x_in <= "01111101"; z_correct<="1101011111110110";
        when 12030 => y_in <= "10101110"; x_in <= "01111110"; z_correct<="1101011110100100";
        when 12031 => y_in <= "10101110"; x_in <= "01111111"; z_correct<="1101011101010010";
        when 12032 => y_in <= "10101111"; x_in <= "10000000"; z_correct<="0010100010000000";
        when 12033 => y_in <= "10101111"; x_in <= "10000001"; z_correct<="0010100000101111";
        when 12034 => y_in <= "10101111"; x_in <= "10000010"; z_correct<="0010011111011110";
        when 12035 => y_in <= "10101111"; x_in <= "10000011"; z_correct<="0010011110001101";
        when 12036 => y_in <= "10101111"; x_in <= "10000100"; z_correct<="0010011100111100";
        when 12037 => y_in <= "10101111"; x_in <= "10000101"; z_correct<="0010011011101011";
        when 12038 => y_in <= "10101111"; x_in <= "10000110"; z_correct<="0010011010011010";
        when 12039 => y_in <= "10101111"; x_in <= "10000111"; z_correct<="0010011001001001";
        when 12040 => y_in <= "10101111"; x_in <= "10001000"; z_correct<="0010010111111000";
        when 12041 => y_in <= "10101111"; x_in <= "10001001"; z_correct<="0010010110100111";
        when 12042 => y_in <= "10101111"; x_in <= "10001010"; z_correct<="0010010101010110";
        when 12043 => y_in <= "10101111"; x_in <= "10001011"; z_correct<="0010010100000101";
        when 12044 => y_in <= "10101111"; x_in <= "10001100"; z_correct<="0010010010110100";
        when 12045 => y_in <= "10101111"; x_in <= "10001101"; z_correct<="0010010001100011";
        when 12046 => y_in <= "10101111"; x_in <= "10001110"; z_correct<="0010010000010010";
        when 12047 => y_in <= "10101111"; x_in <= "10001111"; z_correct<="0010001111000001";
        when 12048 => y_in <= "10101111"; x_in <= "10010000"; z_correct<="0010001101110000";
        when 12049 => y_in <= "10101111"; x_in <= "10010001"; z_correct<="0010001100011111";
        when 12050 => y_in <= "10101111"; x_in <= "10010010"; z_correct<="0010001011001110";
        when 12051 => y_in <= "10101111"; x_in <= "10010011"; z_correct<="0010001001111101";
        when 12052 => y_in <= "10101111"; x_in <= "10010100"; z_correct<="0010001000101100";
        when 12053 => y_in <= "10101111"; x_in <= "10010101"; z_correct<="0010000111011011";
        when 12054 => y_in <= "10101111"; x_in <= "10010110"; z_correct<="0010000110001010";
        when 12055 => y_in <= "10101111"; x_in <= "10010111"; z_correct<="0010000100111001";
        when 12056 => y_in <= "10101111"; x_in <= "10011000"; z_correct<="0010000011101000";
        when 12057 => y_in <= "10101111"; x_in <= "10011001"; z_correct<="0010000010010111";
        when 12058 => y_in <= "10101111"; x_in <= "10011010"; z_correct<="0010000001000110";
        when 12059 => y_in <= "10101111"; x_in <= "10011011"; z_correct<="0001111111110101";
        when 12060 => y_in <= "10101111"; x_in <= "10011100"; z_correct<="0001111110100100";
        when 12061 => y_in <= "10101111"; x_in <= "10011101"; z_correct<="0001111101010011";
        when 12062 => y_in <= "10101111"; x_in <= "10011110"; z_correct<="0001111100000010";
        when 12063 => y_in <= "10101111"; x_in <= "10011111"; z_correct<="0001111010110001";
        when 12064 => y_in <= "10101111"; x_in <= "10100000"; z_correct<="0001111001100000";
        when 12065 => y_in <= "10101111"; x_in <= "10100001"; z_correct<="0001111000001111";
        when 12066 => y_in <= "10101111"; x_in <= "10100010"; z_correct<="0001110110111110";
        when 12067 => y_in <= "10101111"; x_in <= "10100011"; z_correct<="0001110101101101";
        when 12068 => y_in <= "10101111"; x_in <= "10100100"; z_correct<="0001110100011100";
        when 12069 => y_in <= "10101111"; x_in <= "10100101"; z_correct<="0001110011001011";
        when 12070 => y_in <= "10101111"; x_in <= "10100110"; z_correct<="0001110001111010";
        when 12071 => y_in <= "10101111"; x_in <= "10100111"; z_correct<="0001110000101001";
        when 12072 => y_in <= "10101111"; x_in <= "10101000"; z_correct<="0001101111011000";
        when 12073 => y_in <= "10101111"; x_in <= "10101001"; z_correct<="0001101110000111";
        when 12074 => y_in <= "10101111"; x_in <= "10101010"; z_correct<="0001101100110110";
        when 12075 => y_in <= "10101111"; x_in <= "10101011"; z_correct<="0001101011100101";
        when 12076 => y_in <= "10101111"; x_in <= "10101100"; z_correct<="0001101010010100";
        when 12077 => y_in <= "10101111"; x_in <= "10101101"; z_correct<="0001101001000011";
        when 12078 => y_in <= "10101111"; x_in <= "10101110"; z_correct<="0001100111110010";
        when 12079 => y_in <= "10101111"; x_in <= "10101111"; z_correct<="0001100110100001";
        when 12080 => y_in <= "10101111"; x_in <= "10110000"; z_correct<="0001100101010000";
        when 12081 => y_in <= "10101111"; x_in <= "10110001"; z_correct<="0001100011111111";
        when 12082 => y_in <= "10101111"; x_in <= "10110010"; z_correct<="0001100010101110";
        when 12083 => y_in <= "10101111"; x_in <= "10110011"; z_correct<="0001100001011101";
        when 12084 => y_in <= "10101111"; x_in <= "10110100"; z_correct<="0001100000001100";
        when 12085 => y_in <= "10101111"; x_in <= "10110101"; z_correct<="0001011110111011";
        when 12086 => y_in <= "10101111"; x_in <= "10110110"; z_correct<="0001011101101010";
        when 12087 => y_in <= "10101111"; x_in <= "10110111"; z_correct<="0001011100011001";
        when 12088 => y_in <= "10101111"; x_in <= "10111000"; z_correct<="0001011011001000";
        when 12089 => y_in <= "10101111"; x_in <= "10111001"; z_correct<="0001011001110111";
        when 12090 => y_in <= "10101111"; x_in <= "10111010"; z_correct<="0001011000100110";
        when 12091 => y_in <= "10101111"; x_in <= "10111011"; z_correct<="0001010111010101";
        when 12092 => y_in <= "10101111"; x_in <= "10111100"; z_correct<="0001010110000100";
        when 12093 => y_in <= "10101111"; x_in <= "10111101"; z_correct<="0001010100110011";
        when 12094 => y_in <= "10101111"; x_in <= "10111110"; z_correct<="0001010011100010";
        when 12095 => y_in <= "10101111"; x_in <= "10111111"; z_correct<="0001010010010001";
        when 12096 => y_in <= "10101111"; x_in <= "11000000"; z_correct<="0001010001000000";
        when 12097 => y_in <= "10101111"; x_in <= "11000001"; z_correct<="0001001111101111";
        when 12098 => y_in <= "10101111"; x_in <= "11000010"; z_correct<="0001001110011110";
        when 12099 => y_in <= "10101111"; x_in <= "11000011"; z_correct<="0001001101001101";
        when 12100 => y_in <= "10101111"; x_in <= "11000100"; z_correct<="0001001011111100";
        when 12101 => y_in <= "10101111"; x_in <= "11000101"; z_correct<="0001001010101011";
        when 12102 => y_in <= "10101111"; x_in <= "11000110"; z_correct<="0001001001011010";
        when 12103 => y_in <= "10101111"; x_in <= "11000111"; z_correct<="0001001000001001";
        when 12104 => y_in <= "10101111"; x_in <= "11001000"; z_correct<="0001000110111000";
        when 12105 => y_in <= "10101111"; x_in <= "11001001"; z_correct<="0001000101100111";
        when 12106 => y_in <= "10101111"; x_in <= "11001010"; z_correct<="0001000100010110";
        when 12107 => y_in <= "10101111"; x_in <= "11001011"; z_correct<="0001000011000101";
        when 12108 => y_in <= "10101111"; x_in <= "11001100"; z_correct<="0001000001110100";
        when 12109 => y_in <= "10101111"; x_in <= "11001101"; z_correct<="0001000000100011";
        when 12110 => y_in <= "10101111"; x_in <= "11001110"; z_correct<="0000111111010010";
        when 12111 => y_in <= "10101111"; x_in <= "11001111"; z_correct<="0000111110000001";
        when 12112 => y_in <= "10101111"; x_in <= "11010000"; z_correct<="0000111100110000";
        when 12113 => y_in <= "10101111"; x_in <= "11010001"; z_correct<="0000111011011111";
        when 12114 => y_in <= "10101111"; x_in <= "11010010"; z_correct<="0000111010001110";
        when 12115 => y_in <= "10101111"; x_in <= "11010011"; z_correct<="0000111000111101";
        when 12116 => y_in <= "10101111"; x_in <= "11010100"; z_correct<="0000110111101100";
        when 12117 => y_in <= "10101111"; x_in <= "11010101"; z_correct<="0000110110011011";
        when 12118 => y_in <= "10101111"; x_in <= "11010110"; z_correct<="0000110101001010";
        when 12119 => y_in <= "10101111"; x_in <= "11010111"; z_correct<="0000110011111001";
        when 12120 => y_in <= "10101111"; x_in <= "11011000"; z_correct<="0000110010101000";
        when 12121 => y_in <= "10101111"; x_in <= "11011001"; z_correct<="0000110001010111";
        when 12122 => y_in <= "10101111"; x_in <= "11011010"; z_correct<="0000110000000110";
        when 12123 => y_in <= "10101111"; x_in <= "11011011"; z_correct<="0000101110110101";
        when 12124 => y_in <= "10101111"; x_in <= "11011100"; z_correct<="0000101101100100";
        when 12125 => y_in <= "10101111"; x_in <= "11011101"; z_correct<="0000101100010011";
        when 12126 => y_in <= "10101111"; x_in <= "11011110"; z_correct<="0000101011000010";
        when 12127 => y_in <= "10101111"; x_in <= "11011111"; z_correct<="0000101001110001";
        when 12128 => y_in <= "10101111"; x_in <= "11100000"; z_correct<="0000101000100000";
        when 12129 => y_in <= "10101111"; x_in <= "11100001"; z_correct<="0000100111001111";
        when 12130 => y_in <= "10101111"; x_in <= "11100010"; z_correct<="0000100101111110";
        when 12131 => y_in <= "10101111"; x_in <= "11100011"; z_correct<="0000100100101101";
        when 12132 => y_in <= "10101111"; x_in <= "11100100"; z_correct<="0000100011011100";
        when 12133 => y_in <= "10101111"; x_in <= "11100101"; z_correct<="0000100010001011";
        when 12134 => y_in <= "10101111"; x_in <= "11100110"; z_correct<="0000100000111010";
        when 12135 => y_in <= "10101111"; x_in <= "11100111"; z_correct<="0000011111101001";
        when 12136 => y_in <= "10101111"; x_in <= "11101000"; z_correct<="0000011110011000";
        when 12137 => y_in <= "10101111"; x_in <= "11101001"; z_correct<="0000011101000111";
        when 12138 => y_in <= "10101111"; x_in <= "11101010"; z_correct<="0000011011110110";
        when 12139 => y_in <= "10101111"; x_in <= "11101011"; z_correct<="0000011010100101";
        when 12140 => y_in <= "10101111"; x_in <= "11101100"; z_correct<="0000011001010100";
        when 12141 => y_in <= "10101111"; x_in <= "11101101"; z_correct<="0000011000000011";
        when 12142 => y_in <= "10101111"; x_in <= "11101110"; z_correct<="0000010110110010";
        when 12143 => y_in <= "10101111"; x_in <= "11101111"; z_correct<="0000010101100001";
        when 12144 => y_in <= "10101111"; x_in <= "11110000"; z_correct<="0000010100010000";
        when 12145 => y_in <= "10101111"; x_in <= "11110001"; z_correct<="0000010010111111";
        when 12146 => y_in <= "10101111"; x_in <= "11110010"; z_correct<="0000010001101110";
        when 12147 => y_in <= "10101111"; x_in <= "11110011"; z_correct<="0000010000011101";
        when 12148 => y_in <= "10101111"; x_in <= "11110100"; z_correct<="0000001111001100";
        when 12149 => y_in <= "10101111"; x_in <= "11110101"; z_correct<="0000001101111011";
        when 12150 => y_in <= "10101111"; x_in <= "11110110"; z_correct<="0000001100101010";
        when 12151 => y_in <= "10101111"; x_in <= "11110111"; z_correct<="0000001011011001";
        when 12152 => y_in <= "10101111"; x_in <= "11111000"; z_correct<="0000001010001000";
        when 12153 => y_in <= "10101111"; x_in <= "11111001"; z_correct<="0000001000110111";
        when 12154 => y_in <= "10101111"; x_in <= "11111010"; z_correct<="0000000111100110";
        when 12155 => y_in <= "10101111"; x_in <= "11111011"; z_correct<="0000000110010101";
        when 12156 => y_in <= "10101111"; x_in <= "11111100"; z_correct<="0000000101000100";
        when 12157 => y_in <= "10101111"; x_in <= "11111101"; z_correct<="0000000011110011";
        when 12158 => y_in <= "10101111"; x_in <= "11111110"; z_correct<="0000000010100010";
        when 12159 => y_in <= "10101111"; x_in <= "11111111"; z_correct<="0000000001010001";
        when 12160 => y_in <= "10101111"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 12161 => y_in <= "10101111"; x_in <= "00000001"; z_correct<="1111111110101111";
        when 12162 => y_in <= "10101111"; x_in <= "00000010"; z_correct<="1111111101011110";
        when 12163 => y_in <= "10101111"; x_in <= "00000011"; z_correct<="1111111100001101";
        when 12164 => y_in <= "10101111"; x_in <= "00000100"; z_correct<="1111111010111100";
        when 12165 => y_in <= "10101111"; x_in <= "00000101"; z_correct<="1111111001101011";
        when 12166 => y_in <= "10101111"; x_in <= "00000110"; z_correct<="1111111000011010";
        when 12167 => y_in <= "10101111"; x_in <= "00000111"; z_correct<="1111110111001001";
        when 12168 => y_in <= "10101111"; x_in <= "00001000"; z_correct<="1111110101111000";
        when 12169 => y_in <= "10101111"; x_in <= "00001001"; z_correct<="1111110100100111";
        when 12170 => y_in <= "10101111"; x_in <= "00001010"; z_correct<="1111110011010110";
        when 12171 => y_in <= "10101111"; x_in <= "00001011"; z_correct<="1111110010000101";
        when 12172 => y_in <= "10101111"; x_in <= "00001100"; z_correct<="1111110000110100";
        when 12173 => y_in <= "10101111"; x_in <= "00001101"; z_correct<="1111101111100011";
        when 12174 => y_in <= "10101111"; x_in <= "00001110"; z_correct<="1111101110010010";
        when 12175 => y_in <= "10101111"; x_in <= "00001111"; z_correct<="1111101101000001";
        when 12176 => y_in <= "10101111"; x_in <= "00010000"; z_correct<="1111101011110000";
        when 12177 => y_in <= "10101111"; x_in <= "00010001"; z_correct<="1111101010011111";
        when 12178 => y_in <= "10101111"; x_in <= "00010010"; z_correct<="1111101001001110";
        when 12179 => y_in <= "10101111"; x_in <= "00010011"; z_correct<="1111100111111101";
        when 12180 => y_in <= "10101111"; x_in <= "00010100"; z_correct<="1111100110101100";
        when 12181 => y_in <= "10101111"; x_in <= "00010101"; z_correct<="1111100101011011";
        when 12182 => y_in <= "10101111"; x_in <= "00010110"; z_correct<="1111100100001010";
        when 12183 => y_in <= "10101111"; x_in <= "00010111"; z_correct<="1111100010111001";
        when 12184 => y_in <= "10101111"; x_in <= "00011000"; z_correct<="1111100001101000";
        when 12185 => y_in <= "10101111"; x_in <= "00011001"; z_correct<="1111100000010111";
        when 12186 => y_in <= "10101111"; x_in <= "00011010"; z_correct<="1111011111000110";
        when 12187 => y_in <= "10101111"; x_in <= "00011011"; z_correct<="1111011101110101";
        when 12188 => y_in <= "10101111"; x_in <= "00011100"; z_correct<="1111011100100100";
        when 12189 => y_in <= "10101111"; x_in <= "00011101"; z_correct<="1111011011010011";
        when 12190 => y_in <= "10101111"; x_in <= "00011110"; z_correct<="1111011010000010";
        when 12191 => y_in <= "10101111"; x_in <= "00011111"; z_correct<="1111011000110001";
        when 12192 => y_in <= "10101111"; x_in <= "00100000"; z_correct<="1111010111100000";
        when 12193 => y_in <= "10101111"; x_in <= "00100001"; z_correct<="1111010110001111";
        when 12194 => y_in <= "10101111"; x_in <= "00100010"; z_correct<="1111010100111110";
        when 12195 => y_in <= "10101111"; x_in <= "00100011"; z_correct<="1111010011101101";
        when 12196 => y_in <= "10101111"; x_in <= "00100100"; z_correct<="1111010010011100";
        when 12197 => y_in <= "10101111"; x_in <= "00100101"; z_correct<="1111010001001011";
        when 12198 => y_in <= "10101111"; x_in <= "00100110"; z_correct<="1111001111111010";
        when 12199 => y_in <= "10101111"; x_in <= "00100111"; z_correct<="1111001110101001";
        when 12200 => y_in <= "10101111"; x_in <= "00101000"; z_correct<="1111001101011000";
        when 12201 => y_in <= "10101111"; x_in <= "00101001"; z_correct<="1111001100000111";
        when 12202 => y_in <= "10101111"; x_in <= "00101010"; z_correct<="1111001010110110";
        when 12203 => y_in <= "10101111"; x_in <= "00101011"; z_correct<="1111001001100101";
        when 12204 => y_in <= "10101111"; x_in <= "00101100"; z_correct<="1111001000010100";
        when 12205 => y_in <= "10101111"; x_in <= "00101101"; z_correct<="1111000111000011";
        when 12206 => y_in <= "10101111"; x_in <= "00101110"; z_correct<="1111000101110010";
        when 12207 => y_in <= "10101111"; x_in <= "00101111"; z_correct<="1111000100100001";
        when 12208 => y_in <= "10101111"; x_in <= "00110000"; z_correct<="1111000011010000";
        when 12209 => y_in <= "10101111"; x_in <= "00110001"; z_correct<="1111000001111111";
        when 12210 => y_in <= "10101111"; x_in <= "00110010"; z_correct<="1111000000101110";
        when 12211 => y_in <= "10101111"; x_in <= "00110011"; z_correct<="1110111111011101";
        when 12212 => y_in <= "10101111"; x_in <= "00110100"; z_correct<="1110111110001100";
        when 12213 => y_in <= "10101111"; x_in <= "00110101"; z_correct<="1110111100111011";
        when 12214 => y_in <= "10101111"; x_in <= "00110110"; z_correct<="1110111011101010";
        when 12215 => y_in <= "10101111"; x_in <= "00110111"; z_correct<="1110111010011001";
        when 12216 => y_in <= "10101111"; x_in <= "00111000"; z_correct<="1110111001001000";
        when 12217 => y_in <= "10101111"; x_in <= "00111001"; z_correct<="1110110111110111";
        when 12218 => y_in <= "10101111"; x_in <= "00111010"; z_correct<="1110110110100110";
        when 12219 => y_in <= "10101111"; x_in <= "00111011"; z_correct<="1110110101010101";
        when 12220 => y_in <= "10101111"; x_in <= "00111100"; z_correct<="1110110100000100";
        when 12221 => y_in <= "10101111"; x_in <= "00111101"; z_correct<="1110110010110011";
        when 12222 => y_in <= "10101111"; x_in <= "00111110"; z_correct<="1110110001100010";
        when 12223 => y_in <= "10101111"; x_in <= "00111111"; z_correct<="1110110000010001";
        when 12224 => y_in <= "10101111"; x_in <= "01000000"; z_correct<="1110101111000000";
        when 12225 => y_in <= "10101111"; x_in <= "01000001"; z_correct<="1110101101101111";
        when 12226 => y_in <= "10101111"; x_in <= "01000010"; z_correct<="1110101100011110";
        when 12227 => y_in <= "10101111"; x_in <= "01000011"; z_correct<="1110101011001101";
        when 12228 => y_in <= "10101111"; x_in <= "01000100"; z_correct<="1110101001111100";
        when 12229 => y_in <= "10101111"; x_in <= "01000101"; z_correct<="1110101000101011";
        when 12230 => y_in <= "10101111"; x_in <= "01000110"; z_correct<="1110100111011010";
        when 12231 => y_in <= "10101111"; x_in <= "01000111"; z_correct<="1110100110001001";
        when 12232 => y_in <= "10101111"; x_in <= "01001000"; z_correct<="1110100100111000";
        when 12233 => y_in <= "10101111"; x_in <= "01001001"; z_correct<="1110100011100111";
        when 12234 => y_in <= "10101111"; x_in <= "01001010"; z_correct<="1110100010010110";
        when 12235 => y_in <= "10101111"; x_in <= "01001011"; z_correct<="1110100001000101";
        when 12236 => y_in <= "10101111"; x_in <= "01001100"; z_correct<="1110011111110100";
        when 12237 => y_in <= "10101111"; x_in <= "01001101"; z_correct<="1110011110100011";
        when 12238 => y_in <= "10101111"; x_in <= "01001110"; z_correct<="1110011101010010";
        when 12239 => y_in <= "10101111"; x_in <= "01001111"; z_correct<="1110011100000001";
        when 12240 => y_in <= "10101111"; x_in <= "01010000"; z_correct<="1110011010110000";
        when 12241 => y_in <= "10101111"; x_in <= "01010001"; z_correct<="1110011001011111";
        when 12242 => y_in <= "10101111"; x_in <= "01010010"; z_correct<="1110011000001110";
        when 12243 => y_in <= "10101111"; x_in <= "01010011"; z_correct<="1110010110111101";
        when 12244 => y_in <= "10101111"; x_in <= "01010100"; z_correct<="1110010101101100";
        when 12245 => y_in <= "10101111"; x_in <= "01010101"; z_correct<="1110010100011011";
        when 12246 => y_in <= "10101111"; x_in <= "01010110"; z_correct<="1110010011001010";
        when 12247 => y_in <= "10101111"; x_in <= "01010111"; z_correct<="1110010001111001";
        when 12248 => y_in <= "10101111"; x_in <= "01011000"; z_correct<="1110010000101000";
        when 12249 => y_in <= "10101111"; x_in <= "01011001"; z_correct<="1110001111010111";
        when 12250 => y_in <= "10101111"; x_in <= "01011010"; z_correct<="1110001110000110";
        when 12251 => y_in <= "10101111"; x_in <= "01011011"; z_correct<="1110001100110101";
        when 12252 => y_in <= "10101111"; x_in <= "01011100"; z_correct<="1110001011100100";
        when 12253 => y_in <= "10101111"; x_in <= "01011101"; z_correct<="1110001010010011";
        when 12254 => y_in <= "10101111"; x_in <= "01011110"; z_correct<="1110001001000010";
        when 12255 => y_in <= "10101111"; x_in <= "01011111"; z_correct<="1110000111110001";
        when 12256 => y_in <= "10101111"; x_in <= "01100000"; z_correct<="1110000110100000";
        when 12257 => y_in <= "10101111"; x_in <= "01100001"; z_correct<="1110000101001111";
        when 12258 => y_in <= "10101111"; x_in <= "01100010"; z_correct<="1110000011111110";
        when 12259 => y_in <= "10101111"; x_in <= "01100011"; z_correct<="1110000010101101";
        when 12260 => y_in <= "10101111"; x_in <= "01100100"; z_correct<="1110000001011100";
        when 12261 => y_in <= "10101111"; x_in <= "01100101"; z_correct<="1110000000001011";
        when 12262 => y_in <= "10101111"; x_in <= "01100110"; z_correct<="1101111110111010";
        when 12263 => y_in <= "10101111"; x_in <= "01100111"; z_correct<="1101111101101001";
        when 12264 => y_in <= "10101111"; x_in <= "01101000"; z_correct<="1101111100011000";
        when 12265 => y_in <= "10101111"; x_in <= "01101001"; z_correct<="1101111011000111";
        when 12266 => y_in <= "10101111"; x_in <= "01101010"; z_correct<="1101111001110110";
        when 12267 => y_in <= "10101111"; x_in <= "01101011"; z_correct<="1101111000100101";
        when 12268 => y_in <= "10101111"; x_in <= "01101100"; z_correct<="1101110111010100";
        when 12269 => y_in <= "10101111"; x_in <= "01101101"; z_correct<="1101110110000011";
        when 12270 => y_in <= "10101111"; x_in <= "01101110"; z_correct<="1101110100110010";
        when 12271 => y_in <= "10101111"; x_in <= "01101111"; z_correct<="1101110011100001";
        when 12272 => y_in <= "10101111"; x_in <= "01110000"; z_correct<="1101110010010000";
        when 12273 => y_in <= "10101111"; x_in <= "01110001"; z_correct<="1101110000111111";
        when 12274 => y_in <= "10101111"; x_in <= "01110010"; z_correct<="1101101111101110";
        when 12275 => y_in <= "10101111"; x_in <= "01110011"; z_correct<="1101101110011101";
        when 12276 => y_in <= "10101111"; x_in <= "01110100"; z_correct<="1101101101001100";
        when 12277 => y_in <= "10101111"; x_in <= "01110101"; z_correct<="1101101011111011";
        when 12278 => y_in <= "10101111"; x_in <= "01110110"; z_correct<="1101101010101010";
        when 12279 => y_in <= "10101111"; x_in <= "01110111"; z_correct<="1101101001011001";
        when 12280 => y_in <= "10101111"; x_in <= "01111000"; z_correct<="1101101000001000";
        when 12281 => y_in <= "10101111"; x_in <= "01111001"; z_correct<="1101100110110111";
        when 12282 => y_in <= "10101111"; x_in <= "01111010"; z_correct<="1101100101100110";
        when 12283 => y_in <= "10101111"; x_in <= "01111011"; z_correct<="1101100100010101";
        when 12284 => y_in <= "10101111"; x_in <= "01111100"; z_correct<="1101100011000100";
        when 12285 => y_in <= "10101111"; x_in <= "01111101"; z_correct<="1101100001110011";
        when 12286 => y_in <= "10101111"; x_in <= "01111110"; z_correct<="1101100000100010";
        when 12287 => y_in <= "10101111"; x_in <= "01111111"; z_correct<="1101011111010001";
        when 12288 => y_in <= "10110000"; x_in <= "10000000"; z_correct<="0010100000000000";
        when 12289 => y_in <= "10110000"; x_in <= "10000001"; z_correct<="0010011110110000";
        when 12290 => y_in <= "10110000"; x_in <= "10000010"; z_correct<="0010011101100000";
        when 12291 => y_in <= "10110000"; x_in <= "10000011"; z_correct<="0010011100010000";
        when 12292 => y_in <= "10110000"; x_in <= "10000100"; z_correct<="0010011011000000";
        when 12293 => y_in <= "10110000"; x_in <= "10000101"; z_correct<="0010011001110000";
        when 12294 => y_in <= "10110000"; x_in <= "10000110"; z_correct<="0010011000100000";
        when 12295 => y_in <= "10110000"; x_in <= "10000111"; z_correct<="0010010111010000";
        when 12296 => y_in <= "10110000"; x_in <= "10001000"; z_correct<="0010010110000000";
        when 12297 => y_in <= "10110000"; x_in <= "10001001"; z_correct<="0010010100110000";
        when 12298 => y_in <= "10110000"; x_in <= "10001010"; z_correct<="0010010011100000";
        when 12299 => y_in <= "10110000"; x_in <= "10001011"; z_correct<="0010010010010000";
        when 12300 => y_in <= "10110000"; x_in <= "10001100"; z_correct<="0010010001000000";
        when 12301 => y_in <= "10110000"; x_in <= "10001101"; z_correct<="0010001111110000";
        when 12302 => y_in <= "10110000"; x_in <= "10001110"; z_correct<="0010001110100000";
        when 12303 => y_in <= "10110000"; x_in <= "10001111"; z_correct<="0010001101010000";
        when 12304 => y_in <= "10110000"; x_in <= "10010000"; z_correct<="0010001100000000";
        when 12305 => y_in <= "10110000"; x_in <= "10010001"; z_correct<="0010001010110000";
        when 12306 => y_in <= "10110000"; x_in <= "10010010"; z_correct<="0010001001100000";
        when 12307 => y_in <= "10110000"; x_in <= "10010011"; z_correct<="0010001000010000";
        when 12308 => y_in <= "10110000"; x_in <= "10010100"; z_correct<="0010000111000000";
        when 12309 => y_in <= "10110000"; x_in <= "10010101"; z_correct<="0010000101110000";
        when 12310 => y_in <= "10110000"; x_in <= "10010110"; z_correct<="0010000100100000";
        when 12311 => y_in <= "10110000"; x_in <= "10010111"; z_correct<="0010000011010000";
        when 12312 => y_in <= "10110000"; x_in <= "10011000"; z_correct<="0010000010000000";
        when 12313 => y_in <= "10110000"; x_in <= "10011001"; z_correct<="0010000000110000";
        when 12314 => y_in <= "10110000"; x_in <= "10011010"; z_correct<="0001111111100000";
        when 12315 => y_in <= "10110000"; x_in <= "10011011"; z_correct<="0001111110010000";
        when 12316 => y_in <= "10110000"; x_in <= "10011100"; z_correct<="0001111101000000";
        when 12317 => y_in <= "10110000"; x_in <= "10011101"; z_correct<="0001111011110000";
        when 12318 => y_in <= "10110000"; x_in <= "10011110"; z_correct<="0001111010100000";
        when 12319 => y_in <= "10110000"; x_in <= "10011111"; z_correct<="0001111001010000";
        when 12320 => y_in <= "10110000"; x_in <= "10100000"; z_correct<="0001111000000000";
        when 12321 => y_in <= "10110000"; x_in <= "10100001"; z_correct<="0001110110110000";
        when 12322 => y_in <= "10110000"; x_in <= "10100010"; z_correct<="0001110101100000";
        when 12323 => y_in <= "10110000"; x_in <= "10100011"; z_correct<="0001110100010000";
        when 12324 => y_in <= "10110000"; x_in <= "10100100"; z_correct<="0001110011000000";
        when 12325 => y_in <= "10110000"; x_in <= "10100101"; z_correct<="0001110001110000";
        when 12326 => y_in <= "10110000"; x_in <= "10100110"; z_correct<="0001110000100000";
        when 12327 => y_in <= "10110000"; x_in <= "10100111"; z_correct<="0001101111010000";
        when 12328 => y_in <= "10110000"; x_in <= "10101000"; z_correct<="0001101110000000";
        when 12329 => y_in <= "10110000"; x_in <= "10101001"; z_correct<="0001101100110000";
        when 12330 => y_in <= "10110000"; x_in <= "10101010"; z_correct<="0001101011100000";
        when 12331 => y_in <= "10110000"; x_in <= "10101011"; z_correct<="0001101010010000";
        when 12332 => y_in <= "10110000"; x_in <= "10101100"; z_correct<="0001101001000000";
        when 12333 => y_in <= "10110000"; x_in <= "10101101"; z_correct<="0001100111110000";
        when 12334 => y_in <= "10110000"; x_in <= "10101110"; z_correct<="0001100110100000";
        when 12335 => y_in <= "10110000"; x_in <= "10101111"; z_correct<="0001100101010000";
        when 12336 => y_in <= "10110000"; x_in <= "10110000"; z_correct<="0001100100000000";
        when 12337 => y_in <= "10110000"; x_in <= "10110001"; z_correct<="0001100010110000";
        when 12338 => y_in <= "10110000"; x_in <= "10110010"; z_correct<="0001100001100000";
        when 12339 => y_in <= "10110000"; x_in <= "10110011"; z_correct<="0001100000010000";
        when 12340 => y_in <= "10110000"; x_in <= "10110100"; z_correct<="0001011111000000";
        when 12341 => y_in <= "10110000"; x_in <= "10110101"; z_correct<="0001011101110000";
        when 12342 => y_in <= "10110000"; x_in <= "10110110"; z_correct<="0001011100100000";
        when 12343 => y_in <= "10110000"; x_in <= "10110111"; z_correct<="0001011011010000";
        when 12344 => y_in <= "10110000"; x_in <= "10111000"; z_correct<="0001011010000000";
        when 12345 => y_in <= "10110000"; x_in <= "10111001"; z_correct<="0001011000110000";
        when 12346 => y_in <= "10110000"; x_in <= "10111010"; z_correct<="0001010111100000";
        when 12347 => y_in <= "10110000"; x_in <= "10111011"; z_correct<="0001010110010000";
        when 12348 => y_in <= "10110000"; x_in <= "10111100"; z_correct<="0001010101000000";
        when 12349 => y_in <= "10110000"; x_in <= "10111101"; z_correct<="0001010011110000";
        when 12350 => y_in <= "10110000"; x_in <= "10111110"; z_correct<="0001010010100000";
        when 12351 => y_in <= "10110000"; x_in <= "10111111"; z_correct<="0001010001010000";
        when 12352 => y_in <= "10110000"; x_in <= "11000000"; z_correct<="0001010000000000";
        when 12353 => y_in <= "10110000"; x_in <= "11000001"; z_correct<="0001001110110000";
        when 12354 => y_in <= "10110000"; x_in <= "11000010"; z_correct<="0001001101100000";
        when 12355 => y_in <= "10110000"; x_in <= "11000011"; z_correct<="0001001100010000";
        when 12356 => y_in <= "10110000"; x_in <= "11000100"; z_correct<="0001001011000000";
        when 12357 => y_in <= "10110000"; x_in <= "11000101"; z_correct<="0001001001110000";
        when 12358 => y_in <= "10110000"; x_in <= "11000110"; z_correct<="0001001000100000";
        when 12359 => y_in <= "10110000"; x_in <= "11000111"; z_correct<="0001000111010000";
        when 12360 => y_in <= "10110000"; x_in <= "11001000"; z_correct<="0001000110000000";
        when 12361 => y_in <= "10110000"; x_in <= "11001001"; z_correct<="0001000100110000";
        when 12362 => y_in <= "10110000"; x_in <= "11001010"; z_correct<="0001000011100000";
        when 12363 => y_in <= "10110000"; x_in <= "11001011"; z_correct<="0001000010010000";
        when 12364 => y_in <= "10110000"; x_in <= "11001100"; z_correct<="0001000001000000";
        when 12365 => y_in <= "10110000"; x_in <= "11001101"; z_correct<="0000111111110000";
        when 12366 => y_in <= "10110000"; x_in <= "11001110"; z_correct<="0000111110100000";
        when 12367 => y_in <= "10110000"; x_in <= "11001111"; z_correct<="0000111101010000";
        when 12368 => y_in <= "10110000"; x_in <= "11010000"; z_correct<="0000111100000000";
        when 12369 => y_in <= "10110000"; x_in <= "11010001"; z_correct<="0000111010110000";
        when 12370 => y_in <= "10110000"; x_in <= "11010010"; z_correct<="0000111001100000";
        when 12371 => y_in <= "10110000"; x_in <= "11010011"; z_correct<="0000111000010000";
        when 12372 => y_in <= "10110000"; x_in <= "11010100"; z_correct<="0000110111000000";
        when 12373 => y_in <= "10110000"; x_in <= "11010101"; z_correct<="0000110101110000";
        when 12374 => y_in <= "10110000"; x_in <= "11010110"; z_correct<="0000110100100000";
        when 12375 => y_in <= "10110000"; x_in <= "11010111"; z_correct<="0000110011010000";
        when 12376 => y_in <= "10110000"; x_in <= "11011000"; z_correct<="0000110010000000";
        when 12377 => y_in <= "10110000"; x_in <= "11011001"; z_correct<="0000110000110000";
        when 12378 => y_in <= "10110000"; x_in <= "11011010"; z_correct<="0000101111100000";
        when 12379 => y_in <= "10110000"; x_in <= "11011011"; z_correct<="0000101110010000";
        when 12380 => y_in <= "10110000"; x_in <= "11011100"; z_correct<="0000101101000000";
        when 12381 => y_in <= "10110000"; x_in <= "11011101"; z_correct<="0000101011110000";
        when 12382 => y_in <= "10110000"; x_in <= "11011110"; z_correct<="0000101010100000";
        when 12383 => y_in <= "10110000"; x_in <= "11011111"; z_correct<="0000101001010000";
        when 12384 => y_in <= "10110000"; x_in <= "11100000"; z_correct<="0000101000000000";
        when 12385 => y_in <= "10110000"; x_in <= "11100001"; z_correct<="0000100110110000";
        when 12386 => y_in <= "10110000"; x_in <= "11100010"; z_correct<="0000100101100000";
        when 12387 => y_in <= "10110000"; x_in <= "11100011"; z_correct<="0000100100010000";
        when 12388 => y_in <= "10110000"; x_in <= "11100100"; z_correct<="0000100011000000";
        when 12389 => y_in <= "10110000"; x_in <= "11100101"; z_correct<="0000100001110000";
        when 12390 => y_in <= "10110000"; x_in <= "11100110"; z_correct<="0000100000100000";
        when 12391 => y_in <= "10110000"; x_in <= "11100111"; z_correct<="0000011111010000";
        when 12392 => y_in <= "10110000"; x_in <= "11101000"; z_correct<="0000011110000000";
        when 12393 => y_in <= "10110000"; x_in <= "11101001"; z_correct<="0000011100110000";
        when 12394 => y_in <= "10110000"; x_in <= "11101010"; z_correct<="0000011011100000";
        when 12395 => y_in <= "10110000"; x_in <= "11101011"; z_correct<="0000011010010000";
        when 12396 => y_in <= "10110000"; x_in <= "11101100"; z_correct<="0000011001000000";
        when 12397 => y_in <= "10110000"; x_in <= "11101101"; z_correct<="0000010111110000";
        when 12398 => y_in <= "10110000"; x_in <= "11101110"; z_correct<="0000010110100000";
        when 12399 => y_in <= "10110000"; x_in <= "11101111"; z_correct<="0000010101010000";
        when 12400 => y_in <= "10110000"; x_in <= "11110000"; z_correct<="0000010100000000";
        when 12401 => y_in <= "10110000"; x_in <= "11110001"; z_correct<="0000010010110000";
        when 12402 => y_in <= "10110000"; x_in <= "11110010"; z_correct<="0000010001100000";
        when 12403 => y_in <= "10110000"; x_in <= "11110011"; z_correct<="0000010000010000";
        when 12404 => y_in <= "10110000"; x_in <= "11110100"; z_correct<="0000001111000000";
        when 12405 => y_in <= "10110000"; x_in <= "11110101"; z_correct<="0000001101110000";
        when 12406 => y_in <= "10110000"; x_in <= "11110110"; z_correct<="0000001100100000";
        when 12407 => y_in <= "10110000"; x_in <= "11110111"; z_correct<="0000001011010000";
        when 12408 => y_in <= "10110000"; x_in <= "11111000"; z_correct<="0000001010000000";
        when 12409 => y_in <= "10110000"; x_in <= "11111001"; z_correct<="0000001000110000";
        when 12410 => y_in <= "10110000"; x_in <= "11111010"; z_correct<="0000000111100000";
        when 12411 => y_in <= "10110000"; x_in <= "11111011"; z_correct<="0000000110010000";
        when 12412 => y_in <= "10110000"; x_in <= "11111100"; z_correct<="0000000101000000";
        when 12413 => y_in <= "10110000"; x_in <= "11111101"; z_correct<="0000000011110000";
        when 12414 => y_in <= "10110000"; x_in <= "11111110"; z_correct<="0000000010100000";
        when 12415 => y_in <= "10110000"; x_in <= "11111111"; z_correct<="0000000001010000";
        when 12416 => y_in <= "10110000"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 12417 => y_in <= "10110000"; x_in <= "00000001"; z_correct<="1111111110110000";
        when 12418 => y_in <= "10110000"; x_in <= "00000010"; z_correct<="1111111101100000";
        when 12419 => y_in <= "10110000"; x_in <= "00000011"; z_correct<="1111111100010000";
        when 12420 => y_in <= "10110000"; x_in <= "00000100"; z_correct<="1111111011000000";
        when 12421 => y_in <= "10110000"; x_in <= "00000101"; z_correct<="1111111001110000";
        when 12422 => y_in <= "10110000"; x_in <= "00000110"; z_correct<="1111111000100000";
        when 12423 => y_in <= "10110000"; x_in <= "00000111"; z_correct<="1111110111010000";
        when 12424 => y_in <= "10110000"; x_in <= "00001000"; z_correct<="1111110110000000";
        when 12425 => y_in <= "10110000"; x_in <= "00001001"; z_correct<="1111110100110000";
        when 12426 => y_in <= "10110000"; x_in <= "00001010"; z_correct<="1111110011100000";
        when 12427 => y_in <= "10110000"; x_in <= "00001011"; z_correct<="1111110010010000";
        when 12428 => y_in <= "10110000"; x_in <= "00001100"; z_correct<="1111110001000000";
        when 12429 => y_in <= "10110000"; x_in <= "00001101"; z_correct<="1111101111110000";
        when 12430 => y_in <= "10110000"; x_in <= "00001110"; z_correct<="1111101110100000";
        when 12431 => y_in <= "10110000"; x_in <= "00001111"; z_correct<="1111101101010000";
        when 12432 => y_in <= "10110000"; x_in <= "00010000"; z_correct<="1111101100000000";
        when 12433 => y_in <= "10110000"; x_in <= "00010001"; z_correct<="1111101010110000";
        when 12434 => y_in <= "10110000"; x_in <= "00010010"; z_correct<="1111101001100000";
        when 12435 => y_in <= "10110000"; x_in <= "00010011"; z_correct<="1111101000010000";
        when 12436 => y_in <= "10110000"; x_in <= "00010100"; z_correct<="1111100111000000";
        when 12437 => y_in <= "10110000"; x_in <= "00010101"; z_correct<="1111100101110000";
        when 12438 => y_in <= "10110000"; x_in <= "00010110"; z_correct<="1111100100100000";
        when 12439 => y_in <= "10110000"; x_in <= "00010111"; z_correct<="1111100011010000";
        when 12440 => y_in <= "10110000"; x_in <= "00011000"; z_correct<="1111100010000000";
        when 12441 => y_in <= "10110000"; x_in <= "00011001"; z_correct<="1111100000110000";
        when 12442 => y_in <= "10110000"; x_in <= "00011010"; z_correct<="1111011111100000";
        when 12443 => y_in <= "10110000"; x_in <= "00011011"; z_correct<="1111011110010000";
        when 12444 => y_in <= "10110000"; x_in <= "00011100"; z_correct<="1111011101000000";
        when 12445 => y_in <= "10110000"; x_in <= "00011101"; z_correct<="1111011011110000";
        when 12446 => y_in <= "10110000"; x_in <= "00011110"; z_correct<="1111011010100000";
        when 12447 => y_in <= "10110000"; x_in <= "00011111"; z_correct<="1111011001010000";
        when 12448 => y_in <= "10110000"; x_in <= "00100000"; z_correct<="1111011000000000";
        when 12449 => y_in <= "10110000"; x_in <= "00100001"; z_correct<="1111010110110000";
        when 12450 => y_in <= "10110000"; x_in <= "00100010"; z_correct<="1111010101100000";
        when 12451 => y_in <= "10110000"; x_in <= "00100011"; z_correct<="1111010100010000";
        when 12452 => y_in <= "10110000"; x_in <= "00100100"; z_correct<="1111010011000000";
        when 12453 => y_in <= "10110000"; x_in <= "00100101"; z_correct<="1111010001110000";
        when 12454 => y_in <= "10110000"; x_in <= "00100110"; z_correct<="1111010000100000";
        when 12455 => y_in <= "10110000"; x_in <= "00100111"; z_correct<="1111001111010000";
        when 12456 => y_in <= "10110000"; x_in <= "00101000"; z_correct<="1111001110000000";
        when 12457 => y_in <= "10110000"; x_in <= "00101001"; z_correct<="1111001100110000";
        when 12458 => y_in <= "10110000"; x_in <= "00101010"; z_correct<="1111001011100000";
        when 12459 => y_in <= "10110000"; x_in <= "00101011"; z_correct<="1111001010010000";
        when 12460 => y_in <= "10110000"; x_in <= "00101100"; z_correct<="1111001001000000";
        when 12461 => y_in <= "10110000"; x_in <= "00101101"; z_correct<="1111000111110000";
        when 12462 => y_in <= "10110000"; x_in <= "00101110"; z_correct<="1111000110100000";
        when 12463 => y_in <= "10110000"; x_in <= "00101111"; z_correct<="1111000101010000";
        when 12464 => y_in <= "10110000"; x_in <= "00110000"; z_correct<="1111000100000000";
        when 12465 => y_in <= "10110000"; x_in <= "00110001"; z_correct<="1111000010110000";
        when 12466 => y_in <= "10110000"; x_in <= "00110010"; z_correct<="1111000001100000";
        when 12467 => y_in <= "10110000"; x_in <= "00110011"; z_correct<="1111000000010000";
        when 12468 => y_in <= "10110000"; x_in <= "00110100"; z_correct<="1110111111000000";
        when 12469 => y_in <= "10110000"; x_in <= "00110101"; z_correct<="1110111101110000";
        when 12470 => y_in <= "10110000"; x_in <= "00110110"; z_correct<="1110111100100000";
        when 12471 => y_in <= "10110000"; x_in <= "00110111"; z_correct<="1110111011010000";
        when 12472 => y_in <= "10110000"; x_in <= "00111000"; z_correct<="1110111010000000";
        when 12473 => y_in <= "10110000"; x_in <= "00111001"; z_correct<="1110111000110000";
        when 12474 => y_in <= "10110000"; x_in <= "00111010"; z_correct<="1110110111100000";
        when 12475 => y_in <= "10110000"; x_in <= "00111011"; z_correct<="1110110110010000";
        when 12476 => y_in <= "10110000"; x_in <= "00111100"; z_correct<="1110110101000000";
        when 12477 => y_in <= "10110000"; x_in <= "00111101"; z_correct<="1110110011110000";
        when 12478 => y_in <= "10110000"; x_in <= "00111110"; z_correct<="1110110010100000";
        when 12479 => y_in <= "10110000"; x_in <= "00111111"; z_correct<="1110110001010000";
        when 12480 => y_in <= "10110000"; x_in <= "01000000"; z_correct<="1110110000000000";
        when 12481 => y_in <= "10110000"; x_in <= "01000001"; z_correct<="1110101110110000";
        when 12482 => y_in <= "10110000"; x_in <= "01000010"; z_correct<="1110101101100000";
        when 12483 => y_in <= "10110000"; x_in <= "01000011"; z_correct<="1110101100010000";
        when 12484 => y_in <= "10110000"; x_in <= "01000100"; z_correct<="1110101011000000";
        when 12485 => y_in <= "10110000"; x_in <= "01000101"; z_correct<="1110101001110000";
        when 12486 => y_in <= "10110000"; x_in <= "01000110"; z_correct<="1110101000100000";
        when 12487 => y_in <= "10110000"; x_in <= "01000111"; z_correct<="1110100111010000";
        when 12488 => y_in <= "10110000"; x_in <= "01001000"; z_correct<="1110100110000000";
        when 12489 => y_in <= "10110000"; x_in <= "01001001"; z_correct<="1110100100110000";
        when 12490 => y_in <= "10110000"; x_in <= "01001010"; z_correct<="1110100011100000";
        when 12491 => y_in <= "10110000"; x_in <= "01001011"; z_correct<="1110100010010000";
        when 12492 => y_in <= "10110000"; x_in <= "01001100"; z_correct<="1110100001000000";
        when 12493 => y_in <= "10110000"; x_in <= "01001101"; z_correct<="1110011111110000";
        when 12494 => y_in <= "10110000"; x_in <= "01001110"; z_correct<="1110011110100000";
        when 12495 => y_in <= "10110000"; x_in <= "01001111"; z_correct<="1110011101010000";
        when 12496 => y_in <= "10110000"; x_in <= "01010000"; z_correct<="1110011100000000";
        when 12497 => y_in <= "10110000"; x_in <= "01010001"; z_correct<="1110011010110000";
        when 12498 => y_in <= "10110000"; x_in <= "01010010"; z_correct<="1110011001100000";
        when 12499 => y_in <= "10110000"; x_in <= "01010011"; z_correct<="1110011000010000";
        when 12500 => y_in <= "10110000"; x_in <= "01010100"; z_correct<="1110010111000000";
        when 12501 => y_in <= "10110000"; x_in <= "01010101"; z_correct<="1110010101110000";
        when 12502 => y_in <= "10110000"; x_in <= "01010110"; z_correct<="1110010100100000";
        when 12503 => y_in <= "10110000"; x_in <= "01010111"; z_correct<="1110010011010000";
        when 12504 => y_in <= "10110000"; x_in <= "01011000"; z_correct<="1110010010000000";
        when 12505 => y_in <= "10110000"; x_in <= "01011001"; z_correct<="1110010000110000";
        when 12506 => y_in <= "10110000"; x_in <= "01011010"; z_correct<="1110001111100000";
        when 12507 => y_in <= "10110000"; x_in <= "01011011"; z_correct<="1110001110010000";
        when 12508 => y_in <= "10110000"; x_in <= "01011100"; z_correct<="1110001101000000";
        when 12509 => y_in <= "10110000"; x_in <= "01011101"; z_correct<="1110001011110000";
        when 12510 => y_in <= "10110000"; x_in <= "01011110"; z_correct<="1110001010100000";
        when 12511 => y_in <= "10110000"; x_in <= "01011111"; z_correct<="1110001001010000";
        when 12512 => y_in <= "10110000"; x_in <= "01100000"; z_correct<="1110001000000000";
        when 12513 => y_in <= "10110000"; x_in <= "01100001"; z_correct<="1110000110110000";
        when 12514 => y_in <= "10110000"; x_in <= "01100010"; z_correct<="1110000101100000";
        when 12515 => y_in <= "10110000"; x_in <= "01100011"; z_correct<="1110000100010000";
        when 12516 => y_in <= "10110000"; x_in <= "01100100"; z_correct<="1110000011000000";
        when 12517 => y_in <= "10110000"; x_in <= "01100101"; z_correct<="1110000001110000";
        when 12518 => y_in <= "10110000"; x_in <= "01100110"; z_correct<="1110000000100000";
        when 12519 => y_in <= "10110000"; x_in <= "01100111"; z_correct<="1101111111010000";
        when 12520 => y_in <= "10110000"; x_in <= "01101000"; z_correct<="1101111110000000";
        when 12521 => y_in <= "10110000"; x_in <= "01101001"; z_correct<="1101111100110000";
        when 12522 => y_in <= "10110000"; x_in <= "01101010"; z_correct<="1101111011100000";
        when 12523 => y_in <= "10110000"; x_in <= "01101011"; z_correct<="1101111010010000";
        when 12524 => y_in <= "10110000"; x_in <= "01101100"; z_correct<="1101111001000000";
        when 12525 => y_in <= "10110000"; x_in <= "01101101"; z_correct<="1101110111110000";
        when 12526 => y_in <= "10110000"; x_in <= "01101110"; z_correct<="1101110110100000";
        when 12527 => y_in <= "10110000"; x_in <= "01101111"; z_correct<="1101110101010000";
        when 12528 => y_in <= "10110000"; x_in <= "01110000"; z_correct<="1101110100000000";
        when 12529 => y_in <= "10110000"; x_in <= "01110001"; z_correct<="1101110010110000";
        when 12530 => y_in <= "10110000"; x_in <= "01110010"; z_correct<="1101110001100000";
        when 12531 => y_in <= "10110000"; x_in <= "01110011"; z_correct<="1101110000010000";
        when 12532 => y_in <= "10110000"; x_in <= "01110100"; z_correct<="1101101111000000";
        when 12533 => y_in <= "10110000"; x_in <= "01110101"; z_correct<="1101101101110000";
        when 12534 => y_in <= "10110000"; x_in <= "01110110"; z_correct<="1101101100100000";
        when 12535 => y_in <= "10110000"; x_in <= "01110111"; z_correct<="1101101011010000";
        when 12536 => y_in <= "10110000"; x_in <= "01111000"; z_correct<="1101101010000000";
        when 12537 => y_in <= "10110000"; x_in <= "01111001"; z_correct<="1101101000110000";
        when 12538 => y_in <= "10110000"; x_in <= "01111010"; z_correct<="1101100111100000";
        when 12539 => y_in <= "10110000"; x_in <= "01111011"; z_correct<="1101100110010000";
        when 12540 => y_in <= "10110000"; x_in <= "01111100"; z_correct<="1101100101000000";
        when 12541 => y_in <= "10110000"; x_in <= "01111101"; z_correct<="1101100011110000";
        when 12542 => y_in <= "10110000"; x_in <= "01111110"; z_correct<="1101100010100000";
        when 12543 => y_in <= "10110000"; x_in <= "01111111"; z_correct<="1101100001010000";
        when 12544 => y_in <= "10110001"; x_in <= "10000000"; z_correct<="0010011110000000";
        when 12545 => y_in <= "10110001"; x_in <= "10000001"; z_correct<="0010011100110001";
        when 12546 => y_in <= "10110001"; x_in <= "10000010"; z_correct<="0010011011100010";
        when 12547 => y_in <= "10110001"; x_in <= "10000011"; z_correct<="0010011010010011";
        when 12548 => y_in <= "10110001"; x_in <= "10000100"; z_correct<="0010011001000100";
        when 12549 => y_in <= "10110001"; x_in <= "10000101"; z_correct<="0010010111110101";
        when 12550 => y_in <= "10110001"; x_in <= "10000110"; z_correct<="0010010110100110";
        when 12551 => y_in <= "10110001"; x_in <= "10000111"; z_correct<="0010010101010111";
        when 12552 => y_in <= "10110001"; x_in <= "10001000"; z_correct<="0010010100001000";
        when 12553 => y_in <= "10110001"; x_in <= "10001001"; z_correct<="0010010010111001";
        when 12554 => y_in <= "10110001"; x_in <= "10001010"; z_correct<="0010010001101010";
        when 12555 => y_in <= "10110001"; x_in <= "10001011"; z_correct<="0010010000011011";
        when 12556 => y_in <= "10110001"; x_in <= "10001100"; z_correct<="0010001111001100";
        when 12557 => y_in <= "10110001"; x_in <= "10001101"; z_correct<="0010001101111101";
        when 12558 => y_in <= "10110001"; x_in <= "10001110"; z_correct<="0010001100101110";
        when 12559 => y_in <= "10110001"; x_in <= "10001111"; z_correct<="0010001011011111";
        when 12560 => y_in <= "10110001"; x_in <= "10010000"; z_correct<="0010001010010000";
        when 12561 => y_in <= "10110001"; x_in <= "10010001"; z_correct<="0010001001000001";
        when 12562 => y_in <= "10110001"; x_in <= "10010010"; z_correct<="0010000111110010";
        when 12563 => y_in <= "10110001"; x_in <= "10010011"; z_correct<="0010000110100011";
        when 12564 => y_in <= "10110001"; x_in <= "10010100"; z_correct<="0010000101010100";
        when 12565 => y_in <= "10110001"; x_in <= "10010101"; z_correct<="0010000100000101";
        when 12566 => y_in <= "10110001"; x_in <= "10010110"; z_correct<="0010000010110110";
        when 12567 => y_in <= "10110001"; x_in <= "10010111"; z_correct<="0010000001100111";
        when 12568 => y_in <= "10110001"; x_in <= "10011000"; z_correct<="0010000000011000";
        when 12569 => y_in <= "10110001"; x_in <= "10011001"; z_correct<="0001111111001001";
        when 12570 => y_in <= "10110001"; x_in <= "10011010"; z_correct<="0001111101111010";
        when 12571 => y_in <= "10110001"; x_in <= "10011011"; z_correct<="0001111100101011";
        when 12572 => y_in <= "10110001"; x_in <= "10011100"; z_correct<="0001111011011100";
        when 12573 => y_in <= "10110001"; x_in <= "10011101"; z_correct<="0001111010001101";
        when 12574 => y_in <= "10110001"; x_in <= "10011110"; z_correct<="0001111000111110";
        when 12575 => y_in <= "10110001"; x_in <= "10011111"; z_correct<="0001110111101111";
        when 12576 => y_in <= "10110001"; x_in <= "10100000"; z_correct<="0001110110100000";
        when 12577 => y_in <= "10110001"; x_in <= "10100001"; z_correct<="0001110101010001";
        when 12578 => y_in <= "10110001"; x_in <= "10100010"; z_correct<="0001110100000010";
        when 12579 => y_in <= "10110001"; x_in <= "10100011"; z_correct<="0001110010110011";
        when 12580 => y_in <= "10110001"; x_in <= "10100100"; z_correct<="0001110001100100";
        when 12581 => y_in <= "10110001"; x_in <= "10100101"; z_correct<="0001110000010101";
        when 12582 => y_in <= "10110001"; x_in <= "10100110"; z_correct<="0001101111000110";
        when 12583 => y_in <= "10110001"; x_in <= "10100111"; z_correct<="0001101101110111";
        when 12584 => y_in <= "10110001"; x_in <= "10101000"; z_correct<="0001101100101000";
        when 12585 => y_in <= "10110001"; x_in <= "10101001"; z_correct<="0001101011011001";
        when 12586 => y_in <= "10110001"; x_in <= "10101010"; z_correct<="0001101010001010";
        when 12587 => y_in <= "10110001"; x_in <= "10101011"; z_correct<="0001101000111011";
        when 12588 => y_in <= "10110001"; x_in <= "10101100"; z_correct<="0001100111101100";
        when 12589 => y_in <= "10110001"; x_in <= "10101101"; z_correct<="0001100110011101";
        when 12590 => y_in <= "10110001"; x_in <= "10101110"; z_correct<="0001100101001110";
        when 12591 => y_in <= "10110001"; x_in <= "10101111"; z_correct<="0001100011111111";
        when 12592 => y_in <= "10110001"; x_in <= "10110000"; z_correct<="0001100010110000";
        when 12593 => y_in <= "10110001"; x_in <= "10110001"; z_correct<="0001100001100001";
        when 12594 => y_in <= "10110001"; x_in <= "10110010"; z_correct<="0001100000010010";
        when 12595 => y_in <= "10110001"; x_in <= "10110011"; z_correct<="0001011111000011";
        when 12596 => y_in <= "10110001"; x_in <= "10110100"; z_correct<="0001011101110100";
        when 12597 => y_in <= "10110001"; x_in <= "10110101"; z_correct<="0001011100100101";
        when 12598 => y_in <= "10110001"; x_in <= "10110110"; z_correct<="0001011011010110";
        when 12599 => y_in <= "10110001"; x_in <= "10110111"; z_correct<="0001011010000111";
        when 12600 => y_in <= "10110001"; x_in <= "10111000"; z_correct<="0001011000111000";
        when 12601 => y_in <= "10110001"; x_in <= "10111001"; z_correct<="0001010111101001";
        when 12602 => y_in <= "10110001"; x_in <= "10111010"; z_correct<="0001010110011010";
        when 12603 => y_in <= "10110001"; x_in <= "10111011"; z_correct<="0001010101001011";
        when 12604 => y_in <= "10110001"; x_in <= "10111100"; z_correct<="0001010011111100";
        when 12605 => y_in <= "10110001"; x_in <= "10111101"; z_correct<="0001010010101101";
        when 12606 => y_in <= "10110001"; x_in <= "10111110"; z_correct<="0001010001011110";
        when 12607 => y_in <= "10110001"; x_in <= "10111111"; z_correct<="0001010000001111";
        when 12608 => y_in <= "10110001"; x_in <= "11000000"; z_correct<="0001001111000000";
        when 12609 => y_in <= "10110001"; x_in <= "11000001"; z_correct<="0001001101110001";
        when 12610 => y_in <= "10110001"; x_in <= "11000010"; z_correct<="0001001100100010";
        when 12611 => y_in <= "10110001"; x_in <= "11000011"; z_correct<="0001001011010011";
        when 12612 => y_in <= "10110001"; x_in <= "11000100"; z_correct<="0001001010000100";
        when 12613 => y_in <= "10110001"; x_in <= "11000101"; z_correct<="0001001000110101";
        when 12614 => y_in <= "10110001"; x_in <= "11000110"; z_correct<="0001000111100110";
        when 12615 => y_in <= "10110001"; x_in <= "11000111"; z_correct<="0001000110010111";
        when 12616 => y_in <= "10110001"; x_in <= "11001000"; z_correct<="0001000101001000";
        when 12617 => y_in <= "10110001"; x_in <= "11001001"; z_correct<="0001000011111001";
        when 12618 => y_in <= "10110001"; x_in <= "11001010"; z_correct<="0001000010101010";
        when 12619 => y_in <= "10110001"; x_in <= "11001011"; z_correct<="0001000001011011";
        when 12620 => y_in <= "10110001"; x_in <= "11001100"; z_correct<="0001000000001100";
        when 12621 => y_in <= "10110001"; x_in <= "11001101"; z_correct<="0000111110111101";
        when 12622 => y_in <= "10110001"; x_in <= "11001110"; z_correct<="0000111101101110";
        when 12623 => y_in <= "10110001"; x_in <= "11001111"; z_correct<="0000111100011111";
        when 12624 => y_in <= "10110001"; x_in <= "11010000"; z_correct<="0000111011010000";
        when 12625 => y_in <= "10110001"; x_in <= "11010001"; z_correct<="0000111010000001";
        when 12626 => y_in <= "10110001"; x_in <= "11010010"; z_correct<="0000111000110010";
        when 12627 => y_in <= "10110001"; x_in <= "11010011"; z_correct<="0000110111100011";
        when 12628 => y_in <= "10110001"; x_in <= "11010100"; z_correct<="0000110110010100";
        when 12629 => y_in <= "10110001"; x_in <= "11010101"; z_correct<="0000110101000101";
        when 12630 => y_in <= "10110001"; x_in <= "11010110"; z_correct<="0000110011110110";
        when 12631 => y_in <= "10110001"; x_in <= "11010111"; z_correct<="0000110010100111";
        when 12632 => y_in <= "10110001"; x_in <= "11011000"; z_correct<="0000110001011000";
        when 12633 => y_in <= "10110001"; x_in <= "11011001"; z_correct<="0000110000001001";
        when 12634 => y_in <= "10110001"; x_in <= "11011010"; z_correct<="0000101110111010";
        when 12635 => y_in <= "10110001"; x_in <= "11011011"; z_correct<="0000101101101011";
        when 12636 => y_in <= "10110001"; x_in <= "11011100"; z_correct<="0000101100011100";
        when 12637 => y_in <= "10110001"; x_in <= "11011101"; z_correct<="0000101011001101";
        when 12638 => y_in <= "10110001"; x_in <= "11011110"; z_correct<="0000101001111110";
        when 12639 => y_in <= "10110001"; x_in <= "11011111"; z_correct<="0000101000101111";
        when 12640 => y_in <= "10110001"; x_in <= "11100000"; z_correct<="0000100111100000";
        when 12641 => y_in <= "10110001"; x_in <= "11100001"; z_correct<="0000100110010001";
        when 12642 => y_in <= "10110001"; x_in <= "11100010"; z_correct<="0000100101000010";
        when 12643 => y_in <= "10110001"; x_in <= "11100011"; z_correct<="0000100011110011";
        when 12644 => y_in <= "10110001"; x_in <= "11100100"; z_correct<="0000100010100100";
        when 12645 => y_in <= "10110001"; x_in <= "11100101"; z_correct<="0000100001010101";
        when 12646 => y_in <= "10110001"; x_in <= "11100110"; z_correct<="0000100000000110";
        when 12647 => y_in <= "10110001"; x_in <= "11100111"; z_correct<="0000011110110111";
        when 12648 => y_in <= "10110001"; x_in <= "11101000"; z_correct<="0000011101101000";
        when 12649 => y_in <= "10110001"; x_in <= "11101001"; z_correct<="0000011100011001";
        when 12650 => y_in <= "10110001"; x_in <= "11101010"; z_correct<="0000011011001010";
        when 12651 => y_in <= "10110001"; x_in <= "11101011"; z_correct<="0000011001111011";
        when 12652 => y_in <= "10110001"; x_in <= "11101100"; z_correct<="0000011000101100";
        when 12653 => y_in <= "10110001"; x_in <= "11101101"; z_correct<="0000010111011101";
        when 12654 => y_in <= "10110001"; x_in <= "11101110"; z_correct<="0000010110001110";
        when 12655 => y_in <= "10110001"; x_in <= "11101111"; z_correct<="0000010100111111";
        when 12656 => y_in <= "10110001"; x_in <= "11110000"; z_correct<="0000010011110000";
        when 12657 => y_in <= "10110001"; x_in <= "11110001"; z_correct<="0000010010100001";
        when 12658 => y_in <= "10110001"; x_in <= "11110010"; z_correct<="0000010001010010";
        when 12659 => y_in <= "10110001"; x_in <= "11110011"; z_correct<="0000010000000011";
        when 12660 => y_in <= "10110001"; x_in <= "11110100"; z_correct<="0000001110110100";
        when 12661 => y_in <= "10110001"; x_in <= "11110101"; z_correct<="0000001101100101";
        when 12662 => y_in <= "10110001"; x_in <= "11110110"; z_correct<="0000001100010110";
        when 12663 => y_in <= "10110001"; x_in <= "11110111"; z_correct<="0000001011000111";
        when 12664 => y_in <= "10110001"; x_in <= "11111000"; z_correct<="0000001001111000";
        when 12665 => y_in <= "10110001"; x_in <= "11111001"; z_correct<="0000001000101001";
        when 12666 => y_in <= "10110001"; x_in <= "11111010"; z_correct<="0000000111011010";
        when 12667 => y_in <= "10110001"; x_in <= "11111011"; z_correct<="0000000110001011";
        when 12668 => y_in <= "10110001"; x_in <= "11111100"; z_correct<="0000000100111100";
        when 12669 => y_in <= "10110001"; x_in <= "11111101"; z_correct<="0000000011101101";
        when 12670 => y_in <= "10110001"; x_in <= "11111110"; z_correct<="0000000010011110";
        when 12671 => y_in <= "10110001"; x_in <= "11111111"; z_correct<="0000000001001111";
        when 12672 => y_in <= "10110001"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 12673 => y_in <= "10110001"; x_in <= "00000001"; z_correct<="1111111110110001";
        when 12674 => y_in <= "10110001"; x_in <= "00000010"; z_correct<="1111111101100010";
        when 12675 => y_in <= "10110001"; x_in <= "00000011"; z_correct<="1111111100010011";
        when 12676 => y_in <= "10110001"; x_in <= "00000100"; z_correct<="1111111011000100";
        when 12677 => y_in <= "10110001"; x_in <= "00000101"; z_correct<="1111111001110101";
        when 12678 => y_in <= "10110001"; x_in <= "00000110"; z_correct<="1111111000100110";
        when 12679 => y_in <= "10110001"; x_in <= "00000111"; z_correct<="1111110111010111";
        when 12680 => y_in <= "10110001"; x_in <= "00001000"; z_correct<="1111110110001000";
        when 12681 => y_in <= "10110001"; x_in <= "00001001"; z_correct<="1111110100111001";
        when 12682 => y_in <= "10110001"; x_in <= "00001010"; z_correct<="1111110011101010";
        when 12683 => y_in <= "10110001"; x_in <= "00001011"; z_correct<="1111110010011011";
        when 12684 => y_in <= "10110001"; x_in <= "00001100"; z_correct<="1111110001001100";
        when 12685 => y_in <= "10110001"; x_in <= "00001101"; z_correct<="1111101111111101";
        when 12686 => y_in <= "10110001"; x_in <= "00001110"; z_correct<="1111101110101110";
        when 12687 => y_in <= "10110001"; x_in <= "00001111"; z_correct<="1111101101011111";
        when 12688 => y_in <= "10110001"; x_in <= "00010000"; z_correct<="1111101100010000";
        when 12689 => y_in <= "10110001"; x_in <= "00010001"; z_correct<="1111101011000001";
        when 12690 => y_in <= "10110001"; x_in <= "00010010"; z_correct<="1111101001110010";
        when 12691 => y_in <= "10110001"; x_in <= "00010011"; z_correct<="1111101000100011";
        when 12692 => y_in <= "10110001"; x_in <= "00010100"; z_correct<="1111100111010100";
        when 12693 => y_in <= "10110001"; x_in <= "00010101"; z_correct<="1111100110000101";
        when 12694 => y_in <= "10110001"; x_in <= "00010110"; z_correct<="1111100100110110";
        when 12695 => y_in <= "10110001"; x_in <= "00010111"; z_correct<="1111100011100111";
        when 12696 => y_in <= "10110001"; x_in <= "00011000"; z_correct<="1111100010011000";
        when 12697 => y_in <= "10110001"; x_in <= "00011001"; z_correct<="1111100001001001";
        when 12698 => y_in <= "10110001"; x_in <= "00011010"; z_correct<="1111011111111010";
        when 12699 => y_in <= "10110001"; x_in <= "00011011"; z_correct<="1111011110101011";
        when 12700 => y_in <= "10110001"; x_in <= "00011100"; z_correct<="1111011101011100";
        when 12701 => y_in <= "10110001"; x_in <= "00011101"; z_correct<="1111011100001101";
        when 12702 => y_in <= "10110001"; x_in <= "00011110"; z_correct<="1111011010111110";
        when 12703 => y_in <= "10110001"; x_in <= "00011111"; z_correct<="1111011001101111";
        when 12704 => y_in <= "10110001"; x_in <= "00100000"; z_correct<="1111011000100000";
        when 12705 => y_in <= "10110001"; x_in <= "00100001"; z_correct<="1111010111010001";
        when 12706 => y_in <= "10110001"; x_in <= "00100010"; z_correct<="1111010110000010";
        when 12707 => y_in <= "10110001"; x_in <= "00100011"; z_correct<="1111010100110011";
        when 12708 => y_in <= "10110001"; x_in <= "00100100"; z_correct<="1111010011100100";
        when 12709 => y_in <= "10110001"; x_in <= "00100101"; z_correct<="1111010010010101";
        when 12710 => y_in <= "10110001"; x_in <= "00100110"; z_correct<="1111010001000110";
        when 12711 => y_in <= "10110001"; x_in <= "00100111"; z_correct<="1111001111110111";
        when 12712 => y_in <= "10110001"; x_in <= "00101000"; z_correct<="1111001110101000";
        when 12713 => y_in <= "10110001"; x_in <= "00101001"; z_correct<="1111001101011001";
        when 12714 => y_in <= "10110001"; x_in <= "00101010"; z_correct<="1111001100001010";
        when 12715 => y_in <= "10110001"; x_in <= "00101011"; z_correct<="1111001010111011";
        when 12716 => y_in <= "10110001"; x_in <= "00101100"; z_correct<="1111001001101100";
        when 12717 => y_in <= "10110001"; x_in <= "00101101"; z_correct<="1111001000011101";
        when 12718 => y_in <= "10110001"; x_in <= "00101110"; z_correct<="1111000111001110";
        when 12719 => y_in <= "10110001"; x_in <= "00101111"; z_correct<="1111000101111111";
        when 12720 => y_in <= "10110001"; x_in <= "00110000"; z_correct<="1111000100110000";
        when 12721 => y_in <= "10110001"; x_in <= "00110001"; z_correct<="1111000011100001";
        when 12722 => y_in <= "10110001"; x_in <= "00110010"; z_correct<="1111000010010010";
        when 12723 => y_in <= "10110001"; x_in <= "00110011"; z_correct<="1111000001000011";
        when 12724 => y_in <= "10110001"; x_in <= "00110100"; z_correct<="1110111111110100";
        when 12725 => y_in <= "10110001"; x_in <= "00110101"; z_correct<="1110111110100101";
        when 12726 => y_in <= "10110001"; x_in <= "00110110"; z_correct<="1110111101010110";
        when 12727 => y_in <= "10110001"; x_in <= "00110111"; z_correct<="1110111100000111";
        when 12728 => y_in <= "10110001"; x_in <= "00111000"; z_correct<="1110111010111000";
        when 12729 => y_in <= "10110001"; x_in <= "00111001"; z_correct<="1110111001101001";
        when 12730 => y_in <= "10110001"; x_in <= "00111010"; z_correct<="1110111000011010";
        when 12731 => y_in <= "10110001"; x_in <= "00111011"; z_correct<="1110110111001011";
        when 12732 => y_in <= "10110001"; x_in <= "00111100"; z_correct<="1110110101111100";
        when 12733 => y_in <= "10110001"; x_in <= "00111101"; z_correct<="1110110100101101";
        when 12734 => y_in <= "10110001"; x_in <= "00111110"; z_correct<="1110110011011110";
        when 12735 => y_in <= "10110001"; x_in <= "00111111"; z_correct<="1110110010001111";
        when 12736 => y_in <= "10110001"; x_in <= "01000000"; z_correct<="1110110001000000";
        when 12737 => y_in <= "10110001"; x_in <= "01000001"; z_correct<="1110101111110001";
        when 12738 => y_in <= "10110001"; x_in <= "01000010"; z_correct<="1110101110100010";
        when 12739 => y_in <= "10110001"; x_in <= "01000011"; z_correct<="1110101101010011";
        when 12740 => y_in <= "10110001"; x_in <= "01000100"; z_correct<="1110101100000100";
        when 12741 => y_in <= "10110001"; x_in <= "01000101"; z_correct<="1110101010110101";
        when 12742 => y_in <= "10110001"; x_in <= "01000110"; z_correct<="1110101001100110";
        when 12743 => y_in <= "10110001"; x_in <= "01000111"; z_correct<="1110101000010111";
        when 12744 => y_in <= "10110001"; x_in <= "01001000"; z_correct<="1110100111001000";
        when 12745 => y_in <= "10110001"; x_in <= "01001001"; z_correct<="1110100101111001";
        when 12746 => y_in <= "10110001"; x_in <= "01001010"; z_correct<="1110100100101010";
        when 12747 => y_in <= "10110001"; x_in <= "01001011"; z_correct<="1110100011011011";
        when 12748 => y_in <= "10110001"; x_in <= "01001100"; z_correct<="1110100010001100";
        when 12749 => y_in <= "10110001"; x_in <= "01001101"; z_correct<="1110100000111101";
        when 12750 => y_in <= "10110001"; x_in <= "01001110"; z_correct<="1110011111101110";
        when 12751 => y_in <= "10110001"; x_in <= "01001111"; z_correct<="1110011110011111";
        when 12752 => y_in <= "10110001"; x_in <= "01010000"; z_correct<="1110011101010000";
        when 12753 => y_in <= "10110001"; x_in <= "01010001"; z_correct<="1110011100000001";
        when 12754 => y_in <= "10110001"; x_in <= "01010010"; z_correct<="1110011010110010";
        when 12755 => y_in <= "10110001"; x_in <= "01010011"; z_correct<="1110011001100011";
        when 12756 => y_in <= "10110001"; x_in <= "01010100"; z_correct<="1110011000010100";
        when 12757 => y_in <= "10110001"; x_in <= "01010101"; z_correct<="1110010111000101";
        when 12758 => y_in <= "10110001"; x_in <= "01010110"; z_correct<="1110010101110110";
        when 12759 => y_in <= "10110001"; x_in <= "01010111"; z_correct<="1110010100100111";
        when 12760 => y_in <= "10110001"; x_in <= "01011000"; z_correct<="1110010011011000";
        when 12761 => y_in <= "10110001"; x_in <= "01011001"; z_correct<="1110010010001001";
        when 12762 => y_in <= "10110001"; x_in <= "01011010"; z_correct<="1110010000111010";
        when 12763 => y_in <= "10110001"; x_in <= "01011011"; z_correct<="1110001111101011";
        when 12764 => y_in <= "10110001"; x_in <= "01011100"; z_correct<="1110001110011100";
        when 12765 => y_in <= "10110001"; x_in <= "01011101"; z_correct<="1110001101001101";
        when 12766 => y_in <= "10110001"; x_in <= "01011110"; z_correct<="1110001011111110";
        when 12767 => y_in <= "10110001"; x_in <= "01011111"; z_correct<="1110001010101111";
        when 12768 => y_in <= "10110001"; x_in <= "01100000"; z_correct<="1110001001100000";
        when 12769 => y_in <= "10110001"; x_in <= "01100001"; z_correct<="1110001000010001";
        when 12770 => y_in <= "10110001"; x_in <= "01100010"; z_correct<="1110000111000010";
        when 12771 => y_in <= "10110001"; x_in <= "01100011"; z_correct<="1110000101110011";
        when 12772 => y_in <= "10110001"; x_in <= "01100100"; z_correct<="1110000100100100";
        when 12773 => y_in <= "10110001"; x_in <= "01100101"; z_correct<="1110000011010101";
        when 12774 => y_in <= "10110001"; x_in <= "01100110"; z_correct<="1110000010000110";
        when 12775 => y_in <= "10110001"; x_in <= "01100111"; z_correct<="1110000000110111";
        when 12776 => y_in <= "10110001"; x_in <= "01101000"; z_correct<="1101111111101000";
        when 12777 => y_in <= "10110001"; x_in <= "01101001"; z_correct<="1101111110011001";
        when 12778 => y_in <= "10110001"; x_in <= "01101010"; z_correct<="1101111101001010";
        when 12779 => y_in <= "10110001"; x_in <= "01101011"; z_correct<="1101111011111011";
        when 12780 => y_in <= "10110001"; x_in <= "01101100"; z_correct<="1101111010101100";
        when 12781 => y_in <= "10110001"; x_in <= "01101101"; z_correct<="1101111001011101";
        when 12782 => y_in <= "10110001"; x_in <= "01101110"; z_correct<="1101111000001110";
        when 12783 => y_in <= "10110001"; x_in <= "01101111"; z_correct<="1101110110111111";
        when 12784 => y_in <= "10110001"; x_in <= "01110000"; z_correct<="1101110101110000";
        when 12785 => y_in <= "10110001"; x_in <= "01110001"; z_correct<="1101110100100001";
        when 12786 => y_in <= "10110001"; x_in <= "01110010"; z_correct<="1101110011010010";
        when 12787 => y_in <= "10110001"; x_in <= "01110011"; z_correct<="1101110010000011";
        when 12788 => y_in <= "10110001"; x_in <= "01110100"; z_correct<="1101110000110100";
        when 12789 => y_in <= "10110001"; x_in <= "01110101"; z_correct<="1101101111100101";
        when 12790 => y_in <= "10110001"; x_in <= "01110110"; z_correct<="1101101110010110";
        when 12791 => y_in <= "10110001"; x_in <= "01110111"; z_correct<="1101101101000111";
        when 12792 => y_in <= "10110001"; x_in <= "01111000"; z_correct<="1101101011111000";
        when 12793 => y_in <= "10110001"; x_in <= "01111001"; z_correct<="1101101010101001";
        when 12794 => y_in <= "10110001"; x_in <= "01111010"; z_correct<="1101101001011010";
        when 12795 => y_in <= "10110001"; x_in <= "01111011"; z_correct<="1101101000001011";
        when 12796 => y_in <= "10110001"; x_in <= "01111100"; z_correct<="1101100110111100";
        when 12797 => y_in <= "10110001"; x_in <= "01111101"; z_correct<="1101100101101101";
        when 12798 => y_in <= "10110001"; x_in <= "01111110"; z_correct<="1101100100011110";
        when 12799 => y_in <= "10110001"; x_in <= "01111111"; z_correct<="1101100011001111";
        when 12800 => y_in <= "10110010"; x_in <= "10000000"; z_correct<="0010011100000000";
        when 12801 => y_in <= "10110010"; x_in <= "10000001"; z_correct<="0010011010110010";
        when 12802 => y_in <= "10110010"; x_in <= "10000010"; z_correct<="0010011001100100";
        when 12803 => y_in <= "10110010"; x_in <= "10000011"; z_correct<="0010011000010110";
        when 12804 => y_in <= "10110010"; x_in <= "10000100"; z_correct<="0010010111001000";
        when 12805 => y_in <= "10110010"; x_in <= "10000101"; z_correct<="0010010101111010";
        when 12806 => y_in <= "10110010"; x_in <= "10000110"; z_correct<="0010010100101100";
        when 12807 => y_in <= "10110010"; x_in <= "10000111"; z_correct<="0010010011011110";
        when 12808 => y_in <= "10110010"; x_in <= "10001000"; z_correct<="0010010010010000";
        when 12809 => y_in <= "10110010"; x_in <= "10001001"; z_correct<="0010010001000010";
        when 12810 => y_in <= "10110010"; x_in <= "10001010"; z_correct<="0010001111110100";
        when 12811 => y_in <= "10110010"; x_in <= "10001011"; z_correct<="0010001110100110";
        when 12812 => y_in <= "10110010"; x_in <= "10001100"; z_correct<="0010001101011000";
        when 12813 => y_in <= "10110010"; x_in <= "10001101"; z_correct<="0010001100001010";
        when 12814 => y_in <= "10110010"; x_in <= "10001110"; z_correct<="0010001010111100";
        when 12815 => y_in <= "10110010"; x_in <= "10001111"; z_correct<="0010001001101110";
        when 12816 => y_in <= "10110010"; x_in <= "10010000"; z_correct<="0010001000100000";
        when 12817 => y_in <= "10110010"; x_in <= "10010001"; z_correct<="0010000111010010";
        when 12818 => y_in <= "10110010"; x_in <= "10010010"; z_correct<="0010000110000100";
        when 12819 => y_in <= "10110010"; x_in <= "10010011"; z_correct<="0010000100110110";
        when 12820 => y_in <= "10110010"; x_in <= "10010100"; z_correct<="0010000011101000";
        when 12821 => y_in <= "10110010"; x_in <= "10010101"; z_correct<="0010000010011010";
        when 12822 => y_in <= "10110010"; x_in <= "10010110"; z_correct<="0010000001001100";
        when 12823 => y_in <= "10110010"; x_in <= "10010111"; z_correct<="0001111111111110";
        when 12824 => y_in <= "10110010"; x_in <= "10011000"; z_correct<="0001111110110000";
        when 12825 => y_in <= "10110010"; x_in <= "10011001"; z_correct<="0001111101100010";
        when 12826 => y_in <= "10110010"; x_in <= "10011010"; z_correct<="0001111100010100";
        when 12827 => y_in <= "10110010"; x_in <= "10011011"; z_correct<="0001111011000110";
        when 12828 => y_in <= "10110010"; x_in <= "10011100"; z_correct<="0001111001111000";
        when 12829 => y_in <= "10110010"; x_in <= "10011101"; z_correct<="0001111000101010";
        when 12830 => y_in <= "10110010"; x_in <= "10011110"; z_correct<="0001110111011100";
        when 12831 => y_in <= "10110010"; x_in <= "10011111"; z_correct<="0001110110001110";
        when 12832 => y_in <= "10110010"; x_in <= "10100000"; z_correct<="0001110101000000";
        when 12833 => y_in <= "10110010"; x_in <= "10100001"; z_correct<="0001110011110010";
        when 12834 => y_in <= "10110010"; x_in <= "10100010"; z_correct<="0001110010100100";
        when 12835 => y_in <= "10110010"; x_in <= "10100011"; z_correct<="0001110001010110";
        when 12836 => y_in <= "10110010"; x_in <= "10100100"; z_correct<="0001110000001000";
        when 12837 => y_in <= "10110010"; x_in <= "10100101"; z_correct<="0001101110111010";
        when 12838 => y_in <= "10110010"; x_in <= "10100110"; z_correct<="0001101101101100";
        when 12839 => y_in <= "10110010"; x_in <= "10100111"; z_correct<="0001101100011110";
        when 12840 => y_in <= "10110010"; x_in <= "10101000"; z_correct<="0001101011010000";
        when 12841 => y_in <= "10110010"; x_in <= "10101001"; z_correct<="0001101010000010";
        when 12842 => y_in <= "10110010"; x_in <= "10101010"; z_correct<="0001101000110100";
        when 12843 => y_in <= "10110010"; x_in <= "10101011"; z_correct<="0001100111100110";
        when 12844 => y_in <= "10110010"; x_in <= "10101100"; z_correct<="0001100110011000";
        when 12845 => y_in <= "10110010"; x_in <= "10101101"; z_correct<="0001100101001010";
        when 12846 => y_in <= "10110010"; x_in <= "10101110"; z_correct<="0001100011111100";
        when 12847 => y_in <= "10110010"; x_in <= "10101111"; z_correct<="0001100010101110";
        when 12848 => y_in <= "10110010"; x_in <= "10110000"; z_correct<="0001100001100000";
        when 12849 => y_in <= "10110010"; x_in <= "10110001"; z_correct<="0001100000010010";
        when 12850 => y_in <= "10110010"; x_in <= "10110010"; z_correct<="0001011111000100";
        when 12851 => y_in <= "10110010"; x_in <= "10110011"; z_correct<="0001011101110110";
        when 12852 => y_in <= "10110010"; x_in <= "10110100"; z_correct<="0001011100101000";
        when 12853 => y_in <= "10110010"; x_in <= "10110101"; z_correct<="0001011011011010";
        when 12854 => y_in <= "10110010"; x_in <= "10110110"; z_correct<="0001011010001100";
        when 12855 => y_in <= "10110010"; x_in <= "10110111"; z_correct<="0001011000111110";
        when 12856 => y_in <= "10110010"; x_in <= "10111000"; z_correct<="0001010111110000";
        when 12857 => y_in <= "10110010"; x_in <= "10111001"; z_correct<="0001010110100010";
        when 12858 => y_in <= "10110010"; x_in <= "10111010"; z_correct<="0001010101010100";
        when 12859 => y_in <= "10110010"; x_in <= "10111011"; z_correct<="0001010100000110";
        when 12860 => y_in <= "10110010"; x_in <= "10111100"; z_correct<="0001010010111000";
        when 12861 => y_in <= "10110010"; x_in <= "10111101"; z_correct<="0001010001101010";
        when 12862 => y_in <= "10110010"; x_in <= "10111110"; z_correct<="0001010000011100";
        when 12863 => y_in <= "10110010"; x_in <= "10111111"; z_correct<="0001001111001110";
        when 12864 => y_in <= "10110010"; x_in <= "11000000"; z_correct<="0001001110000000";
        when 12865 => y_in <= "10110010"; x_in <= "11000001"; z_correct<="0001001100110010";
        when 12866 => y_in <= "10110010"; x_in <= "11000010"; z_correct<="0001001011100100";
        when 12867 => y_in <= "10110010"; x_in <= "11000011"; z_correct<="0001001010010110";
        when 12868 => y_in <= "10110010"; x_in <= "11000100"; z_correct<="0001001001001000";
        when 12869 => y_in <= "10110010"; x_in <= "11000101"; z_correct<="0001000111111010";
        when 12870 => y_in <= "10110010"; x_in <= "11000110"; z_correct<="0001000110101100";
        when 12871 => y_in <= "10110010"; x_in <= "11000111"; z_correct<="0001000101011110";
        when 12872 => y_in <= "10110010"; x_in <= "11001000"; z_correct<="0001000100010000";
        when 12873 => y_in <= "10110010"; x_in <= "11001001"; z_correct<="0001000011000010";
        when 12874 => y_in <= "10110010"; x_in <= "11001010"; z_correct<="0001000001110100";
        when 12875 => y_in <= "10110010"; x_in <= "11001011"; z_correct<="0001000000100110";
        when 12876 => y_in <= "10110010"; x_in <= "11001100"; z_correct<="0000111111011000";
        when 12877 => y_in <= "10110010"; x_in <= "11001101"; z_correct<="0000111110001010";
        when 12878 => y_in <= "10110010"; x_in <= "11001110"; z_correct<="0000111100111100";
        when 12879 => y_in <= "10110010"; x_in <= "11001111"; z_correct<="0000111011101110";
        when 12880 => y_in <= "10110010"; x_in <= "11010000"; z_correct<="0000111010100000";
        when 12881 => y_in <= "10110010"; x_in <= "11010001"; z_correct<="0000111001010010";
        when 12882 => y_in <= "10110010"; x_in <= "11010010"; z_correct<="0000111000000100";
        when 12883 => y_in <= "10110010"; x_in <= "11010011"; z_correct<="0000110110110110";
        when 12884 => y_in <= "10110010"; x_in <= "11010100"; z_correct<="0000110101101000";
        when 12885 => y_in <= "10110010"; x_in <= "11010101"; z_correct<="0000110100011010";
        when 12886 => y_in <= "10110010"; x_in <= "11010110"; z_correct<="0000110011001100";
        when 12887 => y_in <= "10110010"; x_in <= "11010111"; z_correct<="0000110001111110";
        when 12888 => y_in <= "10110010"; x_in <= "11011000"; z_correct<="0000110000110000";
        when 12889 => y_in <= "10110010"; x_in <= "11011001"; z_correct<="0000101111100010";
        when 12890 => y_in <= "10110010"; x_in <= "11011010"; z_correct<="0000101110010100";
        when 12891 => y_in <= "10110010"; x_in <= "11011011"; z_correct<="0000101101000110";
        when 12892 => y_in <= "10110010"; x_in <= "11011100"; z_correct<="0000101011111000";
        when 12893 => y_in <= "10110010"; x_in <= "11011101"; z_correct<="0000101010101010";
        when 12894 => y_in <= "10110010"; x_in <= "11011110"; z_correct<="0000101001011100";
        when 12895 => y_in <= "10110010"; x_in <= "11011111"; z_correct<="0000101000001110";
        when 12896 => y_in <= "10110010"; x_in <= "11100000"; z_correct<="0000100111000000";
        when 12897 => y_in <= "10110010"; x_in <= "11100001"; z_correct<="0000100101110010";
        when 12898 => y_in <= "10110010"; x_in <= "11100010"; z_correct<="0000100100100100";
        when 12899 => y_in <= "10110010"; x_in <= "11100011"; z_correct<="0000100011010110";
        when 12900 => y_in <= "10110010"; x_in <= "11100100"; z_correct<="0000100010001000";
        when 12901 => y_in <= "10110010"; x_in <= "11100101"; z_correct<="0000100000111010";
        when 12902 => y_in <= "10110010"; x_in <= "11100110"; z_correct<="0000011111101100";
        when 12903 => y_in <= "10110010"; x_in <= "11100111"; z_correct<="0000011110011110";
        when 12904 => y_in <= "10110010"; x_in <= "11101000"; z_correct<="0000011101010000";
        when 12905 => y_in <= "10110010"; x_in <= "11101001"; z_correct<="0000011100000010";
        when 12906 => y_in <= "10110010"; x_in <= "11101010"; z_correct<="0000011010110100";
        when 12907 => y_in <= "10110010"; x_in <= "11101011"; z_correct<="0000011001100110";
        when 12908 => y_in <= "10110010"; x_in <= "11101100"; z_correct<="0000011000011000";
        when 12909 => y_in <= "10110010"; x_in <= "11101101"; z_correct<="0000010111001010";
        when 12910 => y_in <= "10110010"; x_in <= "11101110"; z_correct<="0000010101111100";
        when 12911 => y_in <= "10110010"; x_in <= "11101111"; z_correct<="0000010100101110";
        when 12912 => y_in <= "10110010"; x_in <= "11110000"; z_correct<="0000010011100000";
        when 12913 => y_in <= "10110010"; x_in <= "11110001"; z_correct<="0000010010010010";
        when 12914 => y_in <= "10110010"; x_in <= "11110010"; z_correct<="0000010001000100";
        when 12915 => y_in <= "10110010"; x_in <= "11110011"; z_correct<="0000001111110110";
        when 12916 => y_in <= "10110010"; x_in <= "11110100"; z_correct<="0000001110101000";
        when 12917 => y_in <= "10110010"; x_in <= "11110101"; z_correct<="0000001101011010";
        when 12918 => y_in <= "10110010"; x_in <= "11110110"; z_correct<="0000001100001100";
        when 12919 => y_in <= "10110010"; x_in <= "11110111"; z_correct<="0000001010111110";
        when 12920 => y_in <= "10110010"; x_in <= "11111000"; z_correct<="0000001001110000";
        when 12921 => y_in <= "10110010"; x_in <= "11111001"; z_correct<="0000001000100010";
        when 12922 => y_in <= "10110010"; x_in <= "11111010"; z_correct<="0000000111010100";
        when 12923 => y_in <= "10110010"; x_in <= "11111011"; z_correct<="0000000110000110";
        when 12924 => y_in <= "10110010"; x_in <= "11111100"; z_correct<="0000000100111000";
        when 12925 => y_in <= "10110010"; x_in <= "11111101"; z_correct<="0000000011101010";
        when 12926 => y_in <= "10110010"; x_in <= "11111110"; z_correct<="0000000010011100";
        when 12927 => y_in <= "10110010"; x_in <= "11111111"; z_correct<="0000000001001110";
        when 12928 => y_in <= "10110010"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 12929 => y_in <= "10110010"; x_in <= "00000001"; z_correct<="1111111110110010";
        when 12930 => y_in <= "10110010"; x_in <= "00000010"; z_correct<="1111111101100100";
        when 12931 => y_in <= "10110010"; x_in <= "00000011"; z_correct<="1111111100010110";
        when 12932 => y_in <= "10110010"; x_in <= "00000100"; z_correct<="1111111011001000";
        when 12933 => y_in <= "10110010"; x_in <= "00000101"; z_correct<="1111111001111010";
        when 12934 => y_in <= "10110010"; x_in <= "00000110"; z_correct<="1111111000101100";
        when 12935 => y_in <= "10110010"; x_in <= "00000111"; z_correct<="1111110111011110";
        when 12936 => y_in <= "10110010"; x_in <= "00001000"; z_correct<="1111110110010000";
        when 12937 => y_in <= "10110010"; x_in <= "00001001"; z_correct<="1111110101000010";
        when 12938 => y_in <= "10110010"; x_in <= "00001010"; z_correct<="1111110011110100";
        when 12939 => y_in <= "10110010"; x_in <= "00001011"; z_correct<="1111110010100110";
        when 12940 => y_in <= "10110010"; x_in <= "00001100"; z_correct<="1111110001011000";
        when 12941 => y_in <= "10110010"; x_in <= "00001101"; z_correct<="1111110000001010";
        when 12942 => y_in <= "10110010"; x_in <= "00001110"; z_correct<="1111101110111100";
        when 12943 => y_in <= "10110010"; x_in <= "00001111"; z_correct<="1111101101101110";
        when 12944 => y_in <= "10110010"; x_in <= "00010000"; z_correct<="1111101100100000";
        when 12945 => y_in <= "10110010"; x_in <= "00010001"; z_correct<="1111101011010010";
        when 12946 => y_in <= "10110010"; x_in <= "00010010"; z_correct<="1111101010000100";
        when 12947 => y_in <= "10110010"; x_in <= "00010011"; z_correct<="1111101000110110";
        when 12948 => y_in <= "10110010"; x_in <= "00010100"; z_correct<="1111100111101000";
        when 12949 => y_in <= "10110010"; x_in <= "00010101"; z_correct<="1111100110011010";
        when 12950 => y_in <= "10110010"; x_in <= "00010110"; z_correct<="1111100101001100";
        when 12951 => y_in <= "10110010"; x_in <= "00010111"; z_correct<="1111100011111110";
        when 12952 => y_in <= "10110010"; x_in <= "00011000"; z_correct<="1111100010110000";
        when 12953 => y_in <= "10110010"; x_in <= "00011001"; z_correct<="1111100001100010";
        when 12954 => y_in <= "10110010"; x_in <= "00011010"; z_correct<="1111100000010100";
        when 12955 => y_in <= "10110010"; x_in <= "00011011"; z_correct<="1111011111000110";
        when 12956 => y_in <= "10110010"; x_in <= "00011100"; z_correct<="1111011101111000";
        when 12957 => y_in <= "10110010"; x_in <= "00011101"; z_correct<="1111011100101010";
        when 12958 => y_in <= "10110010"; x_in <= "00011110"; z_correct<="1111011011011100";
        when 12959 => y_in <= "10110010"; x_in <= "00011111"; z_correct<="1111011010001110";
        when 12960 => y_in <= "10110010"; x_in <= "00100000"; z_correct<="1111011001000000";
        when 12961 => y_in <= "10110010"; x_in <= "00100001"; z_correct<="1111010111110010";
        when 12962 => y_in <= "10110010"; x_in <= "00100010"; z_correct<="1111010110100100";
        when 12963 => y_in <= "10110010"; x_in <= "00100011"; z_correct<="1111010101010110";
        when 12964 => y_in <= "10110010"; x_in <= "00100100"; z_correct<="1111010100001000";
        when 12965 => y_in <= "10110010"; x_in <= "00100101"; z_correct<="1111010010111010";
        when 12966 => y_in <= "10110010"; x_in <= "00100110"; z_correct<="1111010001101100";
        when 12967 => y_in <= "10110010"; x_in <= "00100111"; z_correct<="1111010000011110";
        when 12968 => y_in <= "10110010"; x_in <= "00101000"; z_correct<="1111001111010000";
        when 12969 => y_in <= "10110010"; x_in <= "00101001"; z_correct<="1111001110000010";
        when 12970 => y_in <= "10110010"; x_in <= "00101010"; z_correct<="1111001100110100";
        when 12971 => y_in <= "10110010"; x_in <= "00101011"; z_correct<="1111001011100110";
        when 12972 => y_in <= "10110010"; x_in <= "00101100"; z_correct<="1111001010011000";
        when 12973 => y_in <= "10110010"; x_in <= "00101101"; z_correct<="1111001001001010";
        when 12974 => y_in <= "10110010"; x_in <= "00101110"; z_correct<="1111000111111100";
        when 12975 => y_in <= "10110010"; x_in <= "00101111"; z_correct<="1111000110101110";
        when 12976 => y_in <= "10110010"; x_in <= "00110000"; z_correct<="1111000101100000";
        when 12977 => y_in <= "10110010"; x_in <= "00110001"; z_correct<="1111000100010010";
        when 12978 => y_in <= "10110010"; x_in <= "00110010"; z_correct<="1111000011000100";
        when 12979 => y_in <= "10110010"; x_in <= "00110011"; z_correct<="1111000001110110";
        when 12980 => y_in <= "10110010"; x_in <= "00110100"; z_correct<="1111000000101000";
        when 12981 => y_in <= "10110010"; x_in <= "00110101"; z_correct<="1110111111011010";
        when 12982 => y_in <= "10110010"; x_in <= "00110110"; z_correct<="1110111110001100";
        when 12983 => y_in <= "10110010"; x_in <= "00110111"; z_correct<="1110111100111110";
        when 12984 => y_in <= "10110010"; x_in <= "00111000"; z_correct<="1110111011110000";
        when 12985 => y_in <= "10110010"; x_in <= "00111001"; z_correct<="1110111010100010";
        when 12986 => y_in <= "10110010"; x_in <= "00111010"; z_correct<="1110111001010100";
        when 12987 => y_in <= "10110010"; x_in <= "00111011"; z_correct<="1110111000000110";
        when 12988 => y_in <= "10110010"; x_in <= "00111100"; z_correct<="1110110110111000";
        when 12989 => y_in <= "10110010"; x_in <= "00111101"; z_correct<="1110110101101010";
        when 12990 => y_in <= "10110010"; x_in <= "00111110"; z_correct<="1110110100011100";
        when 12991 => y_in <= "10110010"; x_in <= "00111111"; z_correct<="1110110011001110";
        when 12992 => y_in <= "10110010"; x_in <= "01000000"; z_correct<="1110110010000000";
        when 12993 => y_in <= "10110010"; x_in <= "01000001"; z_correct<="1110110000110010";
        when 12994 => y_in <= "10110010"; x_in <= "01000010"; z_correct<="1110101111100100";
        when 12995 => y_in <= "10110010"; x_in <= "01000011"; z_correct<="1110101110010110";
        when 12996 => y_in <= "10110010"; x_in <= "01000100"; z_correct<="1110101101001000";
        when 12997 => y_in <= "10110010"; x_in <= "01000101"; z_correct<="1110101011111010";
        when 12998 => y_in <= "10110010"; x_in <= "01000110"; z_correct<="1110101010101100";
        when 12999 => y_in <= "10110010"; x_in <= "01000111"; z_correct<="1110101001011110";
        when 13000 => y_in <= "10110010"; x_in <= "01001000"; z_correct<="1110101000010000";
        when 13001 => y_in <= "10110010"; x_in <= "01001001"; z_correct<="1110100111000010";
        when 13002 => y_in <= "10110010"; x_in <= "01001010"; z_correct<="1110100101110100";
        when 13003 => y_in <= "10110010"; x_in <= "01001011"; z_correct<="1110100100100110";
        when 13004 => y_in <= "10110010"; x_in <= "01001100"; z_correct<="1110100011011000";
        when 13005 => y_in <= "10110010"; x_in <= "01001101"; z_correct<="1110100010001010";
        when 13006 => y_in <= "10110010"; x_in <= "01001110"; z_correct<="1110100000111100";
        when 13007 => y_in <= "10110010"; x_in <= "01001111"; z_correct<="1110011111101110";
        when 13008 => y_in <= "10110010"; x_in <= "01010000"; z_correct<="1110011110100000";
        when 13009 => y_in <= "10110010"; x_in <= "01010001"; z_correct<="1110011101010010";
        when 13010 => y_in <= "10110010"; x_in <= "01010010"; z_correct<="1110011100000100";
        when 13011 => y_in <= "10110010"; x_in <= "01010011"; z_correct<="1110011010110110";
        when 13012 => y_in <= "10110010"; x_in <= "01010100"; z_correct<="1110011001101000";
        when 13013 => y_in <= "10110010"; x_in <= "01010101"; z_correct<="1110011000011010";
        when 13014 => y_in <= "10110010"; x_in <= "01010110"; z_correct<="1110010111001100";
        when 13015 => y_in <= "10110010"; x_in <= "01010111"; z_correct<="1110010101111110";
        when 13016 => y_in <= "10110010"; x_in <= "01011000"; z_correct<="1110010100110000";
        when 13017 => y_in <= "10110010"; x_in <= "01011001"; z_correct<="1110010011100010";
        when 13018 => y_in <= "10110010"; x_in <= "01011010"; z_correct<="1110010010010100";
        when 13019 => y_in <= "10110010"; x_in <= "01011011"; z_correct<="1110010001000110";
        when 13020 => y_in <= "10110010"; x_in <= "01011100"; z_correct<="1110001111111000";
        when 13021 => y_in <= "10110010"; x_in <= "01011101"; z_correct<="1110001110101010";
        when 13022 => y_in <= "10110010"; x_in <= "01011110"; z_correct<="1110001101011100";
        when 13023 => y_in <= "10110010"; x_in <= "01011111"; z_correct<="1110001100001110";
        when 13024 => y_in <= "10110010"; x_in <= "01100000"; z_correct<="1110001011000000";
        when 13025 => y_in <= "10110010"; x_in <= "01100001"; z_correct<="1110001001110010";
        when 13026 => y_in <= "10110010"; x_in <= "01100010"; z_correct<="1110001000100100";
        when 13027 => y_in <= "10110010"; x_in <= "01100011"; z_correct<="1110000111010110";
        when 13028 => y_in <= "10110010"; x_in <= "01100100"; z_correct<="1110000110001000";
        when 13029 => y_in <= "10110010"; x_in <= "01100101"; z_correct<="1110000100111010";
        when 13030 => y_in <= "10110010"; x_in <= "01100110"; z_correct<="1110000011101100";
        when 13031 => y_in <= "10110010"; x_in <= "01100111"; z_correct<="1110000010011110";
        when 13032 => y_in <= "10110010"; x_in <= "01101000"; z_correct<="1110000001010000";
        when 13033 => y_in <= "10110010"; x_in <= "01101001"; z_correct<="1110000000000010";
        when 13034 => y_in <= "10110010"; x_in <= "01101010"; z_correct<="1101111110110100";
        when 13035 => y_in <= "10110010"; x_in <= "01101011"; z_correct<="1101111101100110";
        when 13036 => y_in <= "10110010"; x_in <= "01101100"; z_correct<="1101111100011000";
        when 13037 => y_in <= "10110010"; x_in <= "01101101"; z_correct<="1101111011001010";
        when 13038 => y_in <= "10110010"; x_in <= "01101110"; z_correct<="1101111001111100";
        when 13039 => y_in <= "10110010"; x_in <= "01101111"; z_correct<="1101111000101110";
        when 13040 => y_in <= "10110010"; x_in <= "01110000"; z_correct<="1101110111100000";
        when 13041 => y_in <= "10110010"; x_in <= "01110001"; z_correct<="1101110110010010";
        when 13042 => y_in <= "10110010"; x_in <= "01110010"; z_correct<="1101110101000100";
        when 13043 => y_in <= "10110010"; x_in <= "01110011"; z_correct<="1101110011110110";
        when 13044 => y_in <= "10110010"; x_in <= "01110100"; z_correct<="1101110010101000";
        when 13045 => y_in <= "10110010"; x_in <= "01110101"; z_correct<="1101110001011010";
        when 13046 => y_in <= "10110010"; x_in <= "01110110"; z_correct<="1101110000001100";
        when 13047 => y_in <= "10110010"; x_in <= "01110111"; z_correct<="1101101110111110";
        when 13048 => y_in <= "10110010"; x_in <= "01111000"; z_correct<="1101101101110000";
        when 13049 => y_in <= "10110010"; x_in <= "01111001"; z_correct<="1101101100100010";
        when 13050 => y_in <= "10110010"; x_in <= "01111010"; z_correct<="1101101011010100";
        when 13051 => y_in <= "10110010"; x_in <= "01111011"; z_correct<="1101101010000110";
        when 13052 => y_in <= "10110010"; x_in <= "01111100"; z_correct<="1101101000111000";
        when 13053 => y_in <= "10110010"; x_in <= "01111101"; z_correct<="1101100111101010";
        when 13054 => y_in <= "10110010"; x_in <= "01111110"; z_correct<="1101100110011100";
        when 13055 => y_in <= "10110010"; x_in <= "01111111"; z_correct<="1101100101001110";
        when 13056 => y_in <= "10110011"; x_in <= "10000000"; z_correct<="0010011010000000";
        when 13057 => y_in <= "10110011"; x_in <= "10000001"; z_correct<="0010011000110011";
        when 13058 => y_in <= "10110011"; x_in <= "10000010"; z_correct<="0010010111100110";
        when 13059 => y_in <= "10110011"; x_in <= "10000011"; z_correct<="0010010110011001";
        when 13060 => y_in <= "10110011"; x_in <= "10000100"; z_correct<="0010010101001100";
        when 13061 => y_in <= "10110011"; x_in <= "10000101"; z_correct<="0010010011111111";
        when 13062 => y_in <= "10110011"; x_in <= "10000110"; z_correct<="0010010010110010";
        when 13063 => y_in <= "10110011"; x_in <= "10000111"; z_correct<="0010010001100101";
        when 13064 => y_in <= "10110011"; x_in <= "10001000"; z_correct<="0010010000011000";
        when 13065 => y_in <= "10110011"; x_in <= "10001001"; z_correct<="0010001111001011";
        when 13066 => y_in <= "10110011"; x_in <= "10001010"; z_correct<="0010001101111110";
        when 13067 => y_in <= "10110011"; x_in <= "10001011"; z_correct<="0010001100110001";
        when 13068 => y_in <= "10110011"; x_in <= "10001100"; z_correct<="0010001011100100";
        when 13069 => y_in <= "10110011"; x_in <= "10001101"; z_correct<="0010001010010111";
        when 13070 => y_in <= "10110011"; x_in <= "10001110"; z_correct<="0010001001001010";
        when 13071 => y_in <= "10110011"; x_in <= "10001111"; z_correct<="0010000111111101";
        when 13072 => y_in <= "10110011"; x_in <= "10010000"; z_correct<="0010000110110000";
        when 13073 => y_in <= "10110011"; x_in <= "10010001"; z_correct<="0010000101100011";
        when 13074 => y_in <= "10110011"; x_in <= "10010010"; z_correct<="0010000100010110";
        when 13075 => y_in <= "10110011"; x_in <= "10010011"; z_correct<="0010000011001001";
        when 13076 => y_in <= "10110011"; x_in <= "10010100"; z_correct<="0010000001111100";
        when 13077 => y_in <= "10110011"; x_in <= "10010101"; z_correct<="0010000000101111";
        when 13078 => y_in <= "10110011"; x_in <= "10010110"; z_correct<="0001111111100010";
        when 13079 => y_in <= "10110011"; x_in <= "10010111"; z_correct<="0001111110010101";
        when 13080 => y_in <= "10110011"; x_in <= "10011000"; z_correct<="0001111101001000";
        when 13081 => y_in <= "10110011"; x_in <= "10011001"; z_correct<="0001111011111011";
        when 13082 => y_in <= "10110011"; x_in <= "10011010"; z_correct<="0001111010101110";
        when 13083 => y_in <= "10110011"; x_in <= "10011011"; z_correct<="0001111001100001";
        when 13084 => y_in <= "10110011"; x_in <= "10011100"; z_correct<="0001111000010100";
        when 13085 => y_in <= "10110011"; x_in <= "10011101"; z_correct<="0001110111000111";
        when 13086 => y_in <= "10110011"; x_in <= "10011110"; z_correct<="0001110101111010";
        when 13087 => y_in <= "10110011"; x_in <= "10011111"; z_correct<="0001110100101101";
        when 13088 => y_in <= "10110011"; x_in <= "10100000"; z_correct<="0001110011100000";
        when 13089 => y_in <= "10110011"; x_in <= "10100001"; z_correct<="0001110010010011";
        when 13090 => y_in <= "10110011"; x_in <= "10100010"; z_correct<="0001110001000110";
        when 13091 => y_in <= "10110011"; x_in <= "10100011"; z_correct<="0001101111111001";
        when 13092 => y_in <= "10110011"; x_in <= "10100100"; z_correct<="0001101110101100";
        when 13093 => y_in <= "10110011"; x_in <= "10100101"; z_correct<="0001101101011111";
        when 13094 => y_in <= "10110011"; x_in <= "10100110"; z_correct<="0001101100010010";
        when 13095 => y_in <= "10110011"; x_in <= "10100111"; z_correct<="0001101011000101";
        when 13096 => y_in <= "10110011"; x_in <= "10101000"; z_correct<="0001101001111000";
        when 13097 => y_in <= "10110011"; x_in <= "10101001"; z_correct<="0001101000101011";
        when 13098 => y_in <= "10110011"; x_in <= "10101010"; z_correct<="0001100111011110";
        when 13099 => y_in <= "10110011"; x_in <= "10101011"; z_correct<="0001100110010001";
        when 13100 => y_in <= "10110011"; x_in <= "10101100"; z_correct<="0001100101000100";
        when 13101 => y_in <= "10110011"; x_in <= "10101101"; z_correct<="0001100011110111";
        when 13102 => y_in <= "10110011"; x_in <= "10101110"; z_correct<="0001100010101010";
        when 13103 => y_in <= "10110011"; x_in <= "10101111"; z_correct<="0001100001011101";
        when 13104 => y_in <= "10110011"; x_in <= "10110000"; z_correct<="0001100000010000";
        when 13105 => y_in <= "10110011"; x_in <= "10110001"; z_correct<="0001011111000011";
        when 13106 => y_in <= "10110011"; x_in <= "10110010"; z_correct<="0001011101110110";
        when 13107 => y_in <= "10110011"; x_in <= "10110011"; z_correct<="0001011100101001";
        when 13108 => y_in <= "10110011"; x_in <= "10110100"; z_correct<="0001011011011100";
        when 13109 => y_in <= "10110011"; x_in <= "10110101"; z_correct<="0001011010001111";
        when 13110 => y_in <= "10110011"; x_in <= "10110110"; z_correct<="0001011001000010";
        when 13111 => y_in <= "10110011"; x_in <= "10110111"; z_correct<="0001010111110101";
        when 13112 => y_in <= "10110011"; x_in <= "10111000"; z_correct<="0001010110101000";
        when 13113 => y_in <= "10110011"; x_in <= "10111001"; z_correct<="0001010101011011";
        when 13114 => y_in <= "10110011"; x_in <= "10111010"; z_correct<="0001010100001110";
        when 13115 => y_in <= "10110011"; x_in <= "10111011"; z_correct<="0001010011000001";
        when 13116 => y_in <= "10110011"; x_in <= "10111100"; z_correct<="0001010001110100";
        when 13117 => y_in <= "10110011"; x_in <= "10111101"; z_correct<="0001010000100111";
        when 13118 => y_in <= "10110011"; x_in <= "10111110"; z_correct<="0001001111011010";
        when 13119 => y_in <= "10110011"; x_in <= "10111111"; z_correct<="0001001110001101";
        when 13120 => y_in <= "10110011"; x_in <= "11000000"; z_correct<="0001001101000000";
        when 13121 => y_in <= "10110011"; x_in <= "11000001"; z_correct<="0001001011110011";
        when 13122 => y_in <= "10110011"; x_in <= "11000010"; z_correct<="0001001010100110";
        when 13123 => y_in <= "10110011"; x_in <= "11000011"; z_correct<="0001001001011001";
        when 13124 => y_in <= "10110011"; x_in <= "11000100"; z_correct<="0001001000001100";
        when 13125 => y_in <= "10110011"; x_in <= "11000101"; z_correct<="0001000110111111";
        when 13126 => y_in <= "10110011"; x_in <= "11000110"; z_correct<="0001000101110010";
        when 13127 => y_in <= "10110011"; x_in <= "11000111"; z_correct<="0001000100100101";
        when 13128 => y_in <= "10110011"; x_in <= "11001000"; z_correct<="0001000011011000";
        when 13129 => y_in <= "10110011"; x_in <= "11001001"; z_correct<="0001000010001011";
        when 13130 => y_in <= "10110011"; x_in <= "11001010"; z_correct<="0001000000111110";
        when 13131 => y_in <= "10110011"; x_in <= "11001011"; z_correct<="0000111111110001";
        when 13132 => y_in <= "10110011"; x_in <= "11001100"; z_correct<="0000111110100100";
        when 13133 => y_in <= "10110011"; x_in <= "11001101"; z_correct<="0000111101010111";
        when 13134 => y_in <= "10110011"; x_in <= "11001110"; z_correct<="0000111100001010";
        when 13135 => y_in <= "10110011"; x_in <= "11001111"; z_correct<="0000111010111101";
        when 13136 => y_in <= "10110011"; x_in <= "11010000"; z_correct<="0000111001110000";
        when 13137 => y_in <= "10110011"; x_in <= "11010001"; z_correct<="0000111000100011";
        when 13138 => y_in <= "10110011"; x_in <= "11010010"; z_correct<="0000110111010110";
        when 13139 => y_in <= "10110011"; x_in <= "11010011"; z_correct<="0000110110001001";
        when 13140 => y_in <= "10110011"; x_in <= "11010100"; z_correct<="0000110100111100";
        when 13141 => y_in <= "10110011"; x_in <= "11010101"; z_correct<="0000110011101111";
        when 13142 => y_in <= "10110011"; x_in <= "11010110"; z_correct<="0000110010100010";
        when 13143 => y_in <= "10110011"; x_in <= "11010111"; z_correct<="0000110001010101";
        when 13144 => y_in <= "10110011"; x_in <= "11011000"; z_correct<="0000110000001000";
        when 13145 => y_in <= "10110011"; x_in <= "11011001"; z_correct<="0000101110111011";
        when 13146 => y_in <= "10110011"; x_in <= "11011010"; z_correct<="0000101101101110";
        when 13147 => y_in <= "10110011"; x_in <= "11011011"; z_correct<="0000101100100001";
        when 13148 => y_in <= "10110011"; x_in <= "11011100"; z_correct<="0000101011010100";
        when 13149 => y_in <= "10110011"; x_in <= "11011101"; z_correct<="0000101010000111";
        when 13150 => y_in <= "10110011"; x_in <= "11011110"; z_correct<="0000101000111010";
        when 13151 => y_in <= "10110011"; x_in <= "11011111"; z_correct<="0000100111101101";
        when 13152 => y_in <= "10110011"; x_in <= "11100000"; z_correct<="0000100110100000";
        when 13153 => y_in <= "10110011"; x_in <= "11100001"; z_correct<="0000100101010011";
        when 13154 => y_in <= "10110011"; x_in <= "11100010"; z_correct<="0000100100000110";
        when 13155 => y_in <= "10110011"; x_in <= "11100011"; z_correct<="0000100010111001";
        when 13156 => y_in <= "10110011"; x_in <= "11100100"; z_correct<="0000100001101100";
        when 13157 => y_in <= "10110011"; x_in <= "11100101"; z_correct<="0000100000011111";
        when 13158 => y_in <= "10110011"; x_in <= "11100110"; z_correct<="0000011111010010";
        when 13159 => y_in <= "10110011"; x_in <= "11100111"; z_correct<="0000011110000101";
        when 13160 => y_in <= "10110011"; x_in <= "11101000"; z_correct<="0000011100111000";
        when 13161 => y_in <= "10110011"; x_in <= "11101001"; z_correct<="0000011011101011";
        when 13162 => y_in <= "10110011"; x_in <= "11101010"; z_correct<="0000011010011110";
        when 13163 => y_in <= "10110011"; x_in <= "11101011"; z_correct<="0000011001010001";
        when 13164 => y_in <= "10110011"; x_in <= "11101100"; z_correct<="0000011000000100";
        when 13165 => y_in <= "10110011"; x_in <= "11101101"; z_correct<="0000010110110111";
        when 13166 => y_in <= "10110011"; x_in <= "11101110"; z_correct<="0000010101101010";
        when 13167 => y_in <= "10110011"; x_in <= "11101111"; z_correct<="0000010100011101";
        when 13168 => y_in <= "10110011"; x_in <= "11110000"; z_correct<="0000010011010000";
        when 13169 => y_in <= "10110011"; x_in <= "11110001"; z_correct<="0000010010000011";
        when 13170 => y_in <= "10110011"; x_in <= "11110010"; z_correct<="0000010000110110";
        when 13171 => y_in <= "10110011"; x_in <= "11110011"; z_correct<="0000001111101001";
        when 13172 => y_in <= "10110011"; x_in <= "11110100"; z_correct<="0000001110011100";
        when 13173 => y_in <= "10110011"; x_in <= "11110101"; z_correct<="0000001101001111";
        when 13174 => y_in <= "10110011"; x_in <= "11110110"; z_correct<="0000001100000010";
        when 13175 => y_in <= "10110011"; x_in <= "11110111"; z_correct<="0000001010110101";
        when 13176 => y_in <= "10110011"; x_in <= "11111000"; z_correct<="0000001001101000";
        when 13177 => y_in <= "10110011"; x_in <= "11111001"; z_correct<="0000001000011011";
        when 13178 => y_in <= "10110011"; x_in <= "11111010"; z_correct<="0000000111001110";
        when 13179 => y_in <= "10110011"; x_in <= "11111011"; z_correct<="0000000110000001";
        when 13180 => y_in <= "10110011"; x_in <= "11111100"; z_correct<="0000000100110100";
        when 13181 => y_in <= "10110011"; x_in <= "11111101"; z_correct<="0000000011100111";
        when 13182 => y_in <= "10110011"; x_in <= "11111110"; z_correct<="0000000010011010";
        when 13183 => y_in <= "10110011"; x_in <= "11111111"; z_correct<="0000000001001101";
        when 13184 => y_in <= "10110011"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 13185 => y_in <= "10110011"; x_in <= "00000001"; z_correct<="1111111110110011";
        when 13186 => y_in <= "10110011"; x_in <= "00000010"; z_correct<="1111111101100110";
        when 13187 => y_in <= "10110011"; x_in <= "00000011"; z_correct<="1111111100011001";
        when 13188 => y_in <= "10110011"; x_in <= "00000100"; z_correct<="1111111011001100";
        when 13189 => y_in <= "10110011"; x_in <= "00000101"; z_correct<="1111111001111111";
        when 13190 => y_in <= "10110011"; x_in <= "00000110"; z_correct<="1111111000110010";
        when 13191 => y_in <= "10110011"; x_in <= "00000111"; z_correct<="1111110111100101";
        when 13192 => y_in <= "10110011"; x_in <= "00001000"; z_correct<="1111110110011000";
        when 13193 => y_in <= "10110011"; x_in <= "00001001"; z_correct<="1111110101001011";
        when 13194 => y_in <= "10110011"; x_in <= "00001010"; z_correct<="1111110011111110";
        when 13195 => y_in <= "10110011"; x_in <= "00001011"; z_correct<="1111110010110001";
        when 13196 => y_in <= "10110011"; x_in <= "00001100"; z_correct<="1111110001100100";
        when 13197 => y_in <= "10110011"; x_in <= "00001101"; z_correct<="1111110000010111";
        when 13198 => y_in <= "10110011"; x_in <= "00001110"; z_correct<="1111101111001010";
        when 13199 => y_in <= "10110011"; x_in <= "00001111"; z_correct<="1111101101111101";
        when 13200 => y_in <= "10110011"; x_in <= "00010000"; z_correct<="1111101100110000";
        when 13201 => y_in <= "10110011"; x_in <= "00010001"; z_correct<="1111101011100011";
        when 13202 => y_in <= "10110011"; x_in <= "00010010"; z_correct<="1111101010010110";
        when 13203 => y_in <= "10110011"; x_in <= "00010011"; z_correct<="1111101001001001";
        when 13204 => y_in <= "10110011"; x_in <= "00010100"; z_correct<="1111100111111100";
        when 13205 => y_in <= "10110011"; x_in <= "00010101"; z_correct<="1111100110101111";
        when 13206 => y_in <= "10110011"; x_in <= "00010110"; z_correct<="1111100101100010";
        when 13207 => y_in <= "10110011"; x_in <= "00010111"; z_correct<="1111100100010101";
        when 13208 => y_in <= "10110011"; x_in <= "00011000"; z_correct<="1111100011001000";
        when 13209 => y_in <= "10110011"; x_in <= "00011001"; z_correct<="1111100001111011";
        when 13210 => y_in <= "10110011"; x_in <= "00011010"; z_correct<="1111100000101110";
        when 13211 => y_in <= "10110011"; x_in <= "00011011"; z_correct<="1111011111100001";
        when 13212 => y_in <= "10110011"; x_in <= "00011100"; z_correct<="1111011110010100";
        when 13213 => y_in <= "10110011"; x_in <= "00011101"; z_correct<="1111011101000111";
        when 13214 => y_in <= "10110011"; x_in <= "00011110"; z_correct<="1111011011111010";
        when 13215 => y_in <= "10110011"; x_in <= "00011111"; z_correct<="1111011010101101";
        when 13216 => y_in <= "10110011"; x_in <= "00100000"; z_correct<="1111011001100000";
        when 13217 => y_in <= "10110011"; x_in <= "00100001"; z_correct<="1111011000010011";
        when 13218 => y_in <= "10110011"; x_in <= "00100010"; z_correct<="1111010111000110";
        when 13219 => y_in <= "10110011"; x_in <= "00100011"; z_correct<="1111010101111001";
        when 13220 => y_in <= "10110011"; x_in <= "00100100"; z_correct<="1111010100101100";
        when 13221 => y_in <= "10110011"; x_in <= "00100101"; z_correct<="1111010011011111";
        when 13222 => y_in <= "10110011"; x_in <= "00100110"; z_correct<="1111010010010010";
        when 13223 => y_in <= "10110011"; x_in <= "00100111"; z_correct<="1111010001000101";
        when 13224 => y_in <= "10110011"; x_in <= "00101000"; z_correct<="1111001111111000";
        when 13225 => y_in <= "10110011"; x_in <= "00101001"; z_correct<="1111001110101011";
        when 13226 => y_in <= "10110011"; x_in <= "00101010"; z_correct<="1111001101011110";
        when 13227 => y_in <= "10110011"; x_in <= "00101011"; z_correct<="1111001100010001";
        when 13228 => y_in <= "10110011"; x_in <= "00101100"; z_correct<="1111001011000100";
        when 13229 => y_in <= "10110011"; x_in <= "00101101"; z_correct<="1111001001110111";
        when 13230 => y_in <= "10110011"; x_in <= "00101110"; z_correct<="1111001000101010";
        when 13231 => y_in <= "10110011"; x_in <= "00101111"; z_correct<="1111000111011101";
        when 13232 => y_in <= "10110011"; x_in <= "00110000"; z_correct<="1111000110010000";
        when 13233 => y_in <= "10110011"; x_in <= "00110001"; z_correct<="1111000101000011";
        when 13234 => y_in <= "10110011"; x_in <= "00110010"; z_correct<="1111000011110110";
        when 13235 => y_in <= "10110011"; x_in <= "00110011"; z_correct<="1111000010101001";
        when 13236 => y_in <= "10110011"; x_in <= "00110100"; z_correct<="1111000001011100";
        when 13237 => y_in <= "10110011"; x_in <= "00110101"; z_correct<="1111000000001111";
        when 13238 => y_in <= "10110011"; x_in <= "00110110"; z_correct<="1110111111000010";
        when 13239 => y_in <= "10110011"; x_in <= "00110111"; z_correct<="1110111101110101";
        when 13240 => y_in <= "10110011"; x_in <= "00111000"; z_correct<="1110111100101000";
        when 13241 => y_in <= "10110011"; x_in <= "00111001"; z_correct<="1110111011011011";
        when 13242 => y_in <= "10110011"; x_in <= "00111010"; z_correct<="1110111010001110";
        when 13243 => y_in <= "10110011"; x_in <= "00111011"; z_correct<="1110111001000001";
        when 13244 => y_in <= "10110011"; x_in <= "00111100"; z_correct<="1110110111110100";
        when 13245 => y_in <= "10110011"; x_in <= "00111101"; z_correct<="1110110110100111";
        when 13246 => y_in <= "10110011"; x_in <= "00111110"; z_correct<="1110110101011010";
        when 13247 => y_in <= "10110011"; x_in <= "00111111"; z_correct<="1110110100001101";
        when 13248 => y_in <= "10110011"; x_in <= "01000000"; z_correct<="1110110011000000";
        when 13249 => y_in <= "10110011"; x_in <= "01000001"; z_correct<="1110110001110011";
        when 13250 => y_in <= "10110011"; x_in <= "01000010"; z_correct<="1110110000100110";
        when 13251 => y_in <= "10110011"; x_in <= "01000011"; z_correct<="1110101111011001";
        when 13252 => y_in <= "10110011"; x_in <= "01000100"; z_correct<="1110101110001100";
        when 13253 => y_in <= "10110011"; x_in <= "01000101"; z_correct<="1110101100111111";
        when 13254 => y_in <= "10110011"; x_in <= "01000110"; z_correct<="1110101011110010";
        when 13255 => y_in <= "10110011"; x_in <= "01000111"; z_correct<="1110101010100101";
        when 13256 => y_in <= "10110011"; x_in <= "01001000"; z_correct<="1110101001011000";
        when 13257 => y_in <= "10110011"; x_in <= "01001001"; z_correct<="1110101000001011";
        when 13258 => y_in <= "10110011"; x_in <= "01001010"; z_correct<="1110100110111110";
        when 13259 => y_in <= "10110011"; x_in <= "01001011"; z_correct<="1110100101110001";
        when 13260 => y_in <= "10110011"; x_in <= "01001100"; z_correct<="1110100100100100";
        when 13261 => y_in <= "10110011"; x_in <= "01001101"; z_correct<="1110100011010111";
        when 13262 => y_in <= "10110011"; x_in <= "01001110"; z_correct<="1110100010001010";
        when 13263 => y_in <= "10110011"; x_in <= "01001111"; z_correct<="1110100000111101";
        when 13264 => y_in <= "10110011"; x_in <= "01010000"; z_correct<="1110011111110000";
        when 13265 => y_in <= "10110011"; x_in <= "01010001"; z_correct<="1110011110100011";
        when 13266 => y_in <= "10110011"; x_in <= "01010010"; z_correct<="1110011101010110";
        when 13267 => y_in <= "10110011"; x_in <= "01010011"; z_correct<="1110011100001001";
        when 13268 => y_in <= "10110011"; x_in <= "01010100"; z_correct<="1110011010111100";
        when 13269 => y_in <= "10110011"; x_in <= "01010101"; z_correct<="1110011001101111";
        when 13270 => y_in <= "10110011"; x_in <= "01010110"; z_correct<="1110011000100010";
        when 13271 => y_in <= "10110011"; x_in <= "01010111"; z_correct<="1110010111010101";
        when 13272 => y_in <= "10110011"; x_in <= "01011000"; z_correct<="1110010110001000";
        when 13273 => y_in <= "10110011"; x_in <= "01011001"; z_correct<="1110010100111011";
        when 13274 => y_in <= "10110011"; x_in <= "01011010"; z_correct<="1110010011101110";
        when 13275 => y_in <= "10110011"; x_in <= "01011011"; z_correct<="1110010010100001";
        when 13276 => y_in <= "10110011"; x_in <= "01011100"; z_correct<="1110010001010100";
        when 13277 => y_in <= "10110011"; x_in <= "01011101"; z_correct<="1110010000000111";
        when 13278 => y_in <= "10110011"; x_in <= "01011110"; z_correct<="1110001110111010";
        when 13279 => y_in <= "10110011"; x_in <= "01011111"; z_correct<="1110001101101101";
        when 13280 => y_in <= "10110011"; x_in <= "01100000"; z_correct<="1110001100100000";
        when 13281 => y_in <= "10110011"; x_in <= "01100001"; z_correct<="1110001011010011";
        when 13282 => y_in <= "10110011"; x_in <= "01100010"; z_correct<="1110001010000110";
        when 13283 => y_in <= "10110011"; x_in <= "01100011"; z_correct<="1110001000111001";
        when 13284 => y_in <= "10110011"; x_in <= "01100100"; z_correct<="1110000111101100";
        when 13285 => y_in <= "10110011"; x_in <= "01100101"; z_correct<="1110000110011111";
        when 13286 => y_in <= "10110011"; x_in <= "01100110"; z_correct<="1110000101010010";
        when 13287 => y_in <= "10110011"; x_in <= "01100111"; z_correct<="1110000100000101";
        when 13288 => y_in <= "10110011"; x_in <= "01101000"; z_correct<="1110000010111000";
        when 13289 => y_in <= "10110011"; x_in <= "01101001"; z_correct<="1110000001101011";
        when 13290 => y_in <= "10110011"; x_in <= "01101010"; z_correct<="1110000000011110";
        when 13291 => y_in <= "10110011"; x_in <= "01101011"; z_correct<="1101111111010001";
        when 13292 => y_in <= "10110011"; x_in <= "01101100"; z_correct<="1101111110000100";
        when 13293 => y_in <= "10110011"; x_in <= "01101101"; z_correct<="1101111100110111";
        when 13294 => y_in <= "10110011"; x_in <= "01101110"; z_correct<="1101111011101010";
        when 13295 => y_in <= "10110011"; x_in <= "01101111"; z_correct<="1101111010011101";
        when 13296 => y_in <= "10110011"; x_in <= "01110000"; z_correct<="1101111001010000";
        when 13297 => y_in <= "10110011"; x_in <= "01110001"; z_correct<="1101111000000011";
        when 13298 => y_in <= "10110011"; x_in <= "01110010"; z_correct<="1101110110110110";
        when 13299 => y_in <= "10110011"; x_in <= "01110011"; z_correct<="1101110101101001";
        when 13300 => y_in <= "10110011"; x_in <= "01110100"; z_correct<="1101110100011100";
        when 13301 => y_in <= "10110011"; x_in <= "01110101"; z_correct<="1101110011001111";
        when 13302 => y_in <= "10110011"; x_in <= "01110110"; z_correct<="1101110010000010";
        when 13303 => y_in <= "10110011"; x_in <= "01110111"; z_correct<="1101110000110101";
        when 13304 => y_in <= "10110011"; x_in <= "01111000"; z_correct<="1101101111101000";
        when 13305 => y_in <= "10110011"; x_in <= "01111001"; z_correct<="1101101110011011";
        when 13306 => y_in <= "10110011"; x_in <= "01111010"; z_correct<="1101101101001110";
        when 13307 => y_in <= "10110011"; x_in <= "01111011"; z_correct<="1101101100000001";
        when 13308 => y_in <= "10110011"; x_in <= "01111100"; z_correct<="1101101010110100";
        when 13309 => y_in <= "10110011"; x_in <= "01111101"; z_correct<="1101101001100111";
        when 13310 => y_in <= "10110011"; x_in <= "01111110"; z_correct<="1101101000011010";
        when 13311 => y_in <= "10110011"; x_in <= "01111111"; z_correct<="1101100111001101";
        when 13312 => y_in <= "10110100"; x_in <= "10000000"; z_correct<="0010011000000000";
        when 13313 => y_in <= "10110100"; x_in <= "10000001"; z_correct<="0010010110110100";
        when 13314 => y_in <= "10110100"; x_in <= "10000010"; z_correct<="0010010101101000";
        when 13315 => y_in <= "10110100"; x_in <= "10000011"; z_correct<="0010010100011100";
        when 13316 => y_in <= "10110100"; x_in <= "10000100"; z_correct<="0010010011010000";
        when 13317 => y_in <= "10110100"; x_in <= "10000101"; z_correct<="0010010010000100";
        when 13318 => y_in <= "10110100"; x_in <= "10000110"; z_correct<="0010010000111000";
        when 13319 => y_in <= "10110100"; x_in <= "10000111"; z_correct<="0010001111101100";
        when 13320 => y_in <= "10110100"; x_in <= "10001000"; z_correct<="0010001110100000";
        when 13321 => y_in <= "10110100"; x_in <= "10001001"; z_correct<="0010001101010100";
        when 13322 => y_in <= "10110100"; x_in <= "10001010"; z_correct<="0010001100001000";
        when 13323 => y_in <= "10110100"; x_in <= "10001011"; z_correct<="0010001010111100";
        when 13324 => y_in <= "10110100"; x_in <= "10001100"; z_correct<="0010001001110000";
        when 13325 => y_in <= "10110100"; x_in <= "10001101"; z_correct<="0010001000100100";
        when 13326 => y_in <= "10110100"; x_in <= "10001110"; z_correct<="0010000111011000";
        when 13327 => y_in <= "10110100"; x_in <= "10001111"; z_correct<="0010000110001100";
        when 13328 => y_in <= "10110100"; x_in <= "10010000"; z_correct<="0010000101000000";
        when 13329 => y_in <= "10110100"; x_in <= "10010001"; z_correct<="0010000011110100";
        when 13330 => y_in <= "10110100"; x_in <= "10010010"; z_correct<="0010000010101000";
        when 13331 => y_in <= "10110100"; x_in <= "10010011"; z_correct<="0010000001011100";
        when 13332 => y_in <= "10110100"; x_in <= "10010100"; z_correct<="0010000000010000";
        when 13333 => y_in <= "10110100"; x_in <= "10010101"; z_correct<="0001111111000100";
        when 13334 => y_in <= "10110100"; x_in <= "10010110"; z_correct<="0001111101111000";
        when 13335 => y_in <= "10110100"; x_in <= "10010111"; z_correct<="0001111100101100";
        when 13336 => y_in <= "10110100"; x_in <= "10011000"; z_correct<="0001111011100000";
        when 13337 => y_in <= "10110100"; x_in <= "10011001"; z_correct<="0001111010010100";
        when 13338 => y_in <= "10110100"; x_in <= "10011010"; z_correct<="0001111001001000";
        when 13339 => y_in <= "10110100"; x_in <= "10011011"; z_correct<="0001110111111100";
        when 13340 => y_in <= "10110100"; x_in <= "10011100"; z_correct<="0001110110110000";
        when 13341 => y_in <= "10110100"; x_in <= "10011101"; z_correct<="0001110101100100";
        when 13342 => y_in <= "10110100"; x_in <= "10011110"; z_correct<="0001110100011000";
        when 13343 => y_in <= "10110100"; x_in <= "10011111"; z_correct<="0001110011001100";
        when 13344 => y_in <= "10110100"; x_in <= "10100000"; z_correct<="0001110010000000";
        when 13345 => y_in <= "10110100"; x_in <= "10100001"; z_correct<="0001110000110100";
        when 13346 => y_in <= "10110100"; x_in <= "10100010"; z_correct<="0001101111101000";
        when 13347 => y_in <= "10110100"; x_in <= "10100011"; z_correct<="0001101110011100";
        when 13348 => y_in <= "10110100"; x_in <= "10100100"; z_correct<="0001101101010000";
        when 13349 => y_in <= "10110100"; x_in <= "10100101"; z_correct<="0001101100000100";
        when 13350 => y_in <= "10110100"; x_in <= "10100110"; z_correct<="0001101010111000";
        when 13351 => y_in <= "10110100"; x_in <= "10100111"; z_correct<="0001101001101100";
        when 13352 => y_in <= "10110100"; x_in <= "10101000"; z_correct<="0001101000100000";
        when 13353 => y_in <= "10110100"; x_in <= "10101001"; z_correct<="0001100111010100";
        when 13354 => y_in <= "10110100"; x_in <= "10101010"; z_correct<="0001100110001000";
        when 13355 => y_in <= "10110100"; x_in <= "10101011"; z_correct<="0001100100111100";
        when 13356 => y_in <= "10110100"; x_in <= "10101100"; z_correct<="0001100011110000";
        when 13357 => y_in <= "10110100"; x_in <= "10101101"; z_correct<="0001100010100100";
        when 13358 => y_in <= "10110100"; x_in <= "10101110"; z_correct<="0001100001011000";
        when 13359 => y_in <= "10110100"; x_in <= "10101111"; z_correct<="0001100000001100";
        when 13360 => y_in <= "10110100"; x_in <= "10110000"; z_correct<="0001011111000000";
        when 13361 => y_in <= "10110100"; x_in <= "10110001"; z_correct<="0001011101110100";
        when 13362 => y_in <= "10110100"; x_in <= "10110010"; z_correct<="0001011100101000";
        when 13363 => y_in <= "10110100"; x_in <= "10110011"; z_correct<="0001011011011100";
        when 13364 => y_in <= "10110100"; x_in <= "10110100"; z_correct<="0001011010010000";
        when 13365 => y_in <= "10110100"; x_in <= "10110101"; z_correct<="0001011001000100";
        when 13366 => y_in <= "10110100"; x_in <= "10110110"; z_correct<="0001010111111000";
        when 13367 => y_in <= "10110100"; x_in <= "10110111"; z_correct<="0001010110101100";
        when 13368 => y_in <= "10110100"; x_in <= "10111000"; z_correct<="0001010101100000";
        when 13369 => y_in <= "10110100"; x_in <= "10111001"; z_correct<="0001010100010100";
        when 13370 => y_in <= "10110100"; x_in <= "10111010"; z_correct<="0001010011001000";
        when 13371 => y_in <= "10110100"; x_in <= "10111011"; z_correct<="0001010001111100";
        when 13372 => y_in <= "10110100"; x_in <= "10111100"; z_correct<="0001010000110000";
        when 13373 => y_in <= "10110100"; x_in <= "10111101"; z_correct<="0001001111100100";
        when 13374 => y_in <= "10110100"; x_in <= "10111110"; z_correct<="0001001110011000";
        when 13375 => y_in <= "10110100"; x_in <= "10111111"; z_correct<="0001001101001100";
        when 13376 => y_in <= "10110100"; x_in <= "11000000"; z_correct<="0001001100000000";
        when 13377 => y_in <= "10110100"; x_in <= "11000001"; z_correct<="0001001010110100";
        when 13378 => y_in <= "10110100"; x_in <= "11000010"; z_correct<="0001001001101000";
        when 13379 => y_in <= "10110100"; x_in <= "11000011"; z_correct<="0001001000011100";
        when 13380 => y_in <= "10110100"; x_in <= "11000100"; z_correct<="0001000111010000";
        when 13381 => y_in <= "10110100"; x_in <= "11000101"; z_correct<="0001000110000100";
        when 13382 => y_in <= "10110100"; x_in <= "11000110"; z_correct<="0001000100111000";
        when 13383 => y_in <= "10110100"; x_in <= "11000111"; z_correct<="0001000011101100";
        when 13384 => y_in <= "10110100"; x_in <= "11001000"; z_correct<="0001000010100000";
        when 13385 => y_in <= "10110100"; x_in <= "11001001"; z_correct<="0001000001010100";
        when 13386 => y_in <= "10110100"; x_in <= "11001010"; z_correct<="0001000000001000";
        when 13387 => y_in <= "10110100"; x_in <= "11001011"; z_correct<="0000111110111100";
        when 13388 => y_in <= "10110100"; x_in <= "11001100"; z_correct<="0000111101110000";
        when 13389 => y_in <= "10110100"; x_in <= "11001101"; z_correct<="0000111100100100";
        when 13390 => y_in <= "10110100"; x_in <= "11001110"; z_correct<="0000111011011000";
        when 13391 => y_in <= "10110100"; x_in <= "11001111"; z_correct<="0000111010001100";
        when 13392 => y_in <= "10110100"; x_in <= "11010000"; z_correct<="0000111001000000";
        when 13393 => y_in <= "10110100"; x_in <= "11010001"; z_correct<="0000110111110100";
        when 13394 => y_in <= "10110100"; x_in <= "11010010"; z_correct<="0000110110101000";
        when 13395 => y_in <= "10110100"; x_in <= "11010011"; z_correct<="0000110101011100";
        when 13396 => y_in <= "10110100"; x_in <= "11010100"; z_correct<="0000110100010000";
        when 13397 => y_in <= "10110100"; x_in <= "11010101"; z_correct<="0000110011000100";
        when 13398 => y_in <= "10110100"; x_in <= "11010110"; z_correct<="0000110001111000";
        when 13399 => y_in <= "10110100"; x_in <= "11010111"; z_correct<="0000110000101100";
        when 13400 => y_in <= "10110100"; x_in <= "11011000"; z_correct<="0000101111100000";
        when 13401 => y_in <= "10110100"; x_in <= "11011001"; z_correct<="0000101110010100";
        when 13402 => y_in <= "10110100"; x_in <= "11011010"; z_correct<="0000101101001000";
        when 13403 => y_in <= "10110100"; x_in <= "11011011"; z_correct<="0000101011111100";
        when 13404 => y_in <= "10110100"; x_in <= "11011100"; z_correct<="0000101010110000";
        when 13405 => y_in <= "10110100"; x_in <= "11011101"; z_correct<="0000101001100100";
        when 13406 => y_in <= "10110100"; x_in <= "11011110"; z_correct<="0000101000011000";
        when 13407 => y_in <= "10110100"; x_in <= "11011111"; z_correct<="0000100111001100";
        when 13408 => y_in <= "10110100"; x_in <= "11100000"; z_correct<="0000100110000000";
        when 13409 => y_in <= "10110100"; x_in <= "11100001"; z_correct<="0000100100110100";
        when 13410 => y_in <= "10110100"; x_in <= "11100010"; z_correct<="0000100011101000";
        when 13411 => y_in <= "10110100"; x_in <= "11100011"; z_correct<="0000100010011100";
        when 13412 => y_in <= "10110100"; x_in <= "11100100"; z_correct<="0000100001010000";
        when 13413 => y_in <= "10110100"; x_in <= "11100101"; z_correct<="0000100000000100";
        when 13414 => y_in <= "10110100"; x_in <= "11100110"; z_correct<="0000011110111000";
        when 13415 => y_in <= "10110100"; x_in <= "11100111"; z_correct<="0000011101101100";
        when 13416 => y_in <= "10110100"; x_in <= "11101000"; z_correct<="0000011100100000";
        when 13417 => y_in <= "10110100"; x_in <= "11101001"; z_correct<="0000011011010100";
        when 13418 => y_in <= "10110100"; x_in <= "11101010"; z_correct<="0000011010001000";
        when 13419 => y_in <= "10110100"; x_in <= "11101011"; z_correct<="0000011000111100";
        when 13420 => y_in <= "10110100"; x_in <= "11101100"; z_correct<="0000010111110000";
        when 13421 => y_in <= "10110100"; x_in <= "11101101"; z_correct<="0000010110100100";
        when 13422 => y_in <= "10110100"; x_in <= "11101110"; z_correct<="0000010101011000";
        when 13423 => y_in <= "10110100"; x_in <= "11101111"; z_correct<="0000010100001100";
        when 13424 => y_in <= "10110100"; x_in <= "11110000"; z_correct<="0000010011000000";
        when 13425 => y_in <= "10110100"; x_in <= "11110001"; z_correct<="0000010001110100";
        when 13426 => y_in <= "10110100"; x_in <= "11110010"; z_correct<="0000010000101000";
        when 13427 => y_in <= "10110100"; x_in <= "11110011"; z_correct<="0000001111011100";
        when 13428 => y_in <= "10110100"; x_in <= "11110100"; z_correct<="0000001110010000";
        when 13429 => y_in <= "10110100"; x_in <= "11110101"; z_correct<="0000001101000100";
        when 13430 => y_in <= "10110100"; x_in <= "11110110"; z_correct<="0000001011111000";
        when 13431 => y_in <= "10110100"; x_in <= "11110111"; z_correct<="0000001010101100";
        when 13432 => y_in <= "10110100"; x_in <= "11111000"; z_correct<="0000001001100000";
        when 13433 => y_in <= "10110100"; x_in <= "11111001"; z_correct<="0000001000010100";
        when 13434 => y_in <= "10110100"; x_in <= "11111010"; z_correct<="0000000111001000";
        when 13435 => y_in <= "10110100"; x_in <= "11111011"; z_correct<="0000000101111100";
        when 13436 => y_in <= "10110100"; x_in <= "11111100"; z_correct<="0000000100110000";
        when 13437 => y_in <= "10110100"; x_in <= "11111101"; z_correct<="0000000011100100";
        when 13438 => y_in <= "10110100"; x_in <= "11111110"; z_correct<="0000000010011000";
        when 13439 => y_in <= "10110100"; x_in <= "11111111"; z_correct<="0000000001001100";
        when 13440 => y_in <= "10110100"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 13441 => y_in <= "10110100"; x_in <= "00000001"; z_correct<="1111111110110100";
        when 13442 => y_in <= "10110100"; x_in <= "00000010"; z_correct<="1111111101101000";
        when 13443 => y_in <= "10110100"; x_in <= "00000011"; z_correct<="1111111100011100";
        when 13444 => y_in <= "10110100"; x_in <= "00000100"; z_correct<="1111111011010000";
        when 13445 => y_in <= "10110100"; x_in <= "00000101"; z_correct<="1111111010000100";
        when 13446 => y_in <= "10110100"; x_in <= "00000110"; z_correct<="1111111000111000";
        when 13447 => y_in <= "10110100"; x_in <= "00000111"; z_correct<="1111110111101100";
        when 13448 => y_in <= "10110100"; x_in <= "00001000"; z_correct<="1111110110100000";
        when 13449 => y_in <= "10110100"; x_in <= "00001001"; z_correct<="1111110101010100";
        when 13450 => y_in <= "10110100"; x_in <= "00001010"; z_correct<="1111110100001000";
        when 13451 => y_in <= "10110100"; x_in <= "00001011"; z_correct<="1111110010111100";
        when 13452 => y_in <= "10110100"; x_in <= "00001100"; z_correct<="1111110001110000";
        when 13453 => y_in <= "10110100"; x_in <= "00001101"; z_correct<="1111110000100100";
        when 13454 => y_in <= "10110100"; x_in <= "00001110"; z_correct<="1111101111011000";
        when 13455 => y_in <= "10110100"; x_in <= "00001111"; z_correct<="1111101110001100";
        when 13456 => y_in <= "10110100"; x_in <= "00010000"; z_correct<="1111101101000000";
        when 13457 => y_in <= "10110100"; x_in <= "00010001"; z_correct<="1111101011110100";
        when 13458 => y_in <= "10110100"; x_in <= "00010010"; z_correct<="1111101010101000";
        when 13459 => y_in <= "10110100"; x_in <= "00010011"; z_correct<="1111101001011100";
        when 13460 => y_in <= "10110100"; x_in <= "00010100"; z_correct<="1111101000010000";
        when 13461 => y_in <= "10110100"; x_in <= "00010101"; z_correct<="1111100111000100";
        when 13462 => y_in <= "10110100"; x_in <= "00010110"; z_correct<="1111100101111000";
        when 13463 => y_in <= "10110100"; x_in <= "00010111"; z_correct<="1111100100101100";
        when 13464 => y_in <= "10110100"; x_in <= "00011000"; z_correct<="1111100011100000";
        when 13465 => y_in <= "10110100"; x_in <= "00011001"; z_correct<="1111100010010100";
        when 13466 => y_in <= "10110100"; x_in <= "00011010"; z_correct<="1111100001001000";
        when 13467 => y_in <= "10110100"; x_in <= "00011011"; z_correct<="1111011111111100";
        when 13468 => y_in <= "10110100"; x_in <= "00011100"; z_correct<="1111011110110000";
        when 13469 => y_in <= "10110100"; x_in <= "00011101"; z_correct<="1111011101100100";
        when 13470 => y_in <= "10110100"; x_in <= "00011110"; z_correct<="1111011100011000";
        when 13471 => y_in <= "10110100"; x_in <= "00011111"; z_correct<="1111011011001100";
        when 13472 => y_in <= "10110100"; x_in <= "00100000"; z_correct<="1111011010000000";
        when 13473 => y_in <= "10110100"; x_in <= "00100001"; z_correct<="1111011000110100";
        when 13474 => y_in <= "10110100"; x_in <= "00100010"; z_correct<="1111010111101000";
        when 13475 => y_in <= "10110100"; x_in <= "00100011"; z_correct<="1111010110011100";
        when 13476 => y_in <= "10110100"; x_in <= "00100100"; z_correct<="1111010101010000";
        when 13477 => y_in <= "10110100"; x_in <= "00100101"; z_correct<="1111010100000100";
        when 13478 => y_in <= "10110100"; x_in <= "00100110"; z_correct<="1111010010111000";
        when 13479 => y_in <= "10110100"; x_in <= "00100111"; z_correct<="1111010001101100";
        when 13480 => y_in <= "10110100"; x_in <= "00101000"; z_correct<="1111010000100000";
        when 13481 => y_in <= "10110100"; x_in <= "00101001"; z_correct<="1111001111010100";
        when 13482 => y_in <= "10110100"; x_in <= "00101010"; z_correct<="1111001110001000";
        when 13483 => y_in <= "10110100"; x_in <= "00101011"; z_correct<="1111001100111100";
        when 13484 => y_in <= "10110100"; x_in <= "00101100"; z_correct<="1111001011110000";
        when 13485 => y_in <= "10110100"; x_in <= "00101101"; z_correct<="1111001010100100";
        when 13486 => y_in <= "10110100"; x_in <= "00101110"; z_correct<="1111001001011000";
        when 13487 => y_in <= "10110100"; x_in <= "00101111"; z_correct<="1111001000001100";
        when 13488 => y_in <= "10110100"; x_in <= "00110000"; z_correct<="1111000111000000";
        when 13489 => y_in <= "10110100"; x_in <= "00110001"; z_correct<="1111000101110100";
        when 13490 => y_in <= "10110100"; x_in <= "00110010"; z_correct<="1111000100101000";
        when 13491 => y_in <= "10110100"; x_in <= "00110011"; z_correct<="1111000011011100";
        when 13492 => y_in <= "10110100"; x_in <= "00110100"; z_correct<="1111000010010000";
        when 13493 => y_in <= "10110100"; x_in <= "00110101"; z_correct<="1111000001000100";
        when 13494 => y_in <= "10110100"; x_in <= "00110110"; z_correct<="1110111111111000";
        when 13495 => y_in <= "10110100"; x_in <= "00110111"; z_correct<="1110111110101100";
        when 13496 => y_in <= "10110100"; x_in <= "00111000"; z_correct<="1110111101100000";
        when 13497 => y_in <= "10110100"; x_in <= "00111001"; z_correct<="1110111100010100";
        when 13498 => y_in <= "10110100"; x_in <= "00111010"; z_correct<="1110111011001000";
        when 13499 => y_in <= "10110100"; x_in <= "00111011"; z_correct<="1110111001111100";
        when 13500 => y_in <= "10110100"; x_in <= "00111100"; z_correct<="1110111000110000";
        when 13501 => y_in <= "10110100"; x_in <= "00111101"; z_correct<="1110110111100100";
        when 13502 => y_in <= "10110100"; x_in <= "00111110"; z_correct<="1110110110011000";
        when 13503 => y_in <= "10110100"; x_in <= "00111111"; z_correct<="1110110101001100";
        when 13504 => y_in <= "10110100"; x_in <= "01000000"; z_correct<="1110110100000000";
        when 13505 => y_in <= "10110100"; x_in <= "01000001"; z_correct<="1110110010110100";
        when 13506 => y_in <= "10110100"; x_in <= "01000010"; z_correct<="1110110001101000";
        when 13507 => y_in <= "10110100"; x_in <= "01000011"; z_correct<="1110110000011100";
        when 13508 => y_in <= "10110100"; x_in <= "01000100"; z_correct<="1110101111010000";
        when 13509 => y_in <= "10110100"; x_in <= "01000101"; z_correct<="1110101110000100";
        when 13510 => y_in <= "10110100"; x_in <= "01000110"; z_correct<="1110101100111000";
        when 13511 => y_in <= "10110100"; x_in <= "01000111"; z_correct<="1110101011101100";
        when 13512 => y_in <= "10110100"; x_in <= "01001000"; z_correct<="1110101010100000";
        when 13513 => y_in <= "10110100"; x_in <= "01001001"; z_correct<="1110101001010100";
        when 13514 => y_in <= "10110100"; x_in <= "01001010"; z_correct<="1110101000001000";
        when 13515 => y_in <= "10110100"; x_in <= "01001011"; z_correct<="1110100110111100";
        when 13516 => y_in <= "10110100"; x_in <= "01001100"; z_correct<="1110100101110000";
        when 13517 => y_in <= "10110100"; x_in <= "01001101"; z_correct<="1110100100100100";
        when 13518 => y_in <= "10110100"; x_in <= "01001110"; z_correct<="1110100011011000";
        when 13519 => y_in <= "10110100"; x_in <= "01001111"; z_correct<="1110100010001100";
        when 13520 => y_in <= "10110100"; x_in <= "01010000"; z_correct<="1110100001000000";
        when 13521 => y_in <= "10110100"; x_in <= "01010001"; z_correct<="1110011111110100";
        when 13522 => y_in <= "10110100"; x_in <= "01010010"; z_correct<="1110011110101000";
        when 13523 => y_in <= "10110100"; x_in <= "01010011"; z_correct<="1110011101011100";
        when 13524 => y_in <= "10110100"; x_in <= "01010100"; z_correct<="1110011100010000";
        when 13525 => y_in <= "10110100"; x_in <= "01010101"; z_correct<="1110011011000100";
        when 13526 => y_in <= "10110100"; x_in <= "01010110"; z_correct<="1110011001111000";
        when 13527 => y_in <= "10110100"; x_in <= "01010111"; z_correct<="1110011000101100";
        when 13528 => y_in <= "10110100"; x_in <= "01011000"; z_correct<="1110010111100000";
        when 13529 => y_in <= "10110100"; x_in <= "01011001"; z_correct<="1110010110010100";
        when 13530 => y_in <= "10110100"; x_in <= "01011010"; z_correct<="1110010101001000";
        when 13531 => y_in <= "10110100"; x_in <= "01011011"; z_correct<="1110010011111100";
        when 13532 => y_in <= "10110100"; x_in <= "01011100"; z_correct<="1110010010110000";
        when 13533 => y_in <= "10110100"; x_in <= "01011101"; z_correct<="1110010001100100";
        when 13534 => y_in <= "10110100"; x_in <= "01011110"; z_correct<="1110010000011000";
        when 13535 => y_in <= "10110100"; x_in <= "01011111"; z_correct<="1110001111001100";
        when 13536 => y_in <= "10110100"; x_in <= "01100000"; z_correct<="1110001110000000";
        when 13537 => y_in <= "10110100"; x_in <= "01100001"; z_correct<="1110001100110100";
        when 13538 => y_in <= "10110100"; x_in <= "01100010"; z_correct<="1110001011101000";
        when 13539 => y_in <= "10110100"; x_in <= "01100011"; z_correct<="1110001010011100";
        when 13540 => y_in <= "10110100"; x_in <= "01100100"; z_correct<="1110001001010000";
        when 13541 => y_in <= "10110100"; x_in <= "01100101"; z_correct<="1110001000000100";
        when 13542 => y_in <= "10110100"; x_in <= "01100110"; z_correct<="1110000110111000";
        when 13543 => y_in <= "10110100"; x_in <= "01100111"; z_correct<="1110000101101100";
        when 13544 => y_in <= "10110100"; x_in <= "01101000"; z_correct<="1110000100100000";
        when 13545 => y_in <= "10110100"; x_in <= "01101001"; z_correct<="1110000011010100";
        when 13546 => y_in <= "10110100"; x_in <= "01101010"; z_correct<="1110000010001000";
        when 13547 => y_in <= "10110100"; x_in <= "01101011"; z_correct<="1110000000111100";
        when 13548 => y_in <= "10110100"; x_in <= "01101100"; z_correct<="1101111111110000";
        when 13549 => y_in <= "10110100"; x_in <= "01101101"; z_correct<="1101111110100100";
        when 13550 => y_in <= "10110100"; x_in <= "01101110"; z_correct<="1101111101011000";
        when 13551 => y_in <= "10110100"; x_in <= "01101111"; z_correct<="1101111100001100";
        when 13552 => y_in <= "10110100"; x_in <= "01110000"; z_correct<="1101111011000000";
        when 13553 => y_in <= "10110100"; x_in <= "01110001"; z_correct<="1101111001110100";
        when 13554 => y_in <= "10110100"; x_in <= "01110010"; z_correct<="1101111000101000";
        when 13555 => y_in <= "10110100"; x_in <= "01110011"; z_correct<="1101110111011100";
        when 13556 => y_in <= "10110100"; x_in <= "01110100"; z_correct<="1101110110010000";
        when 13557 => y_in <= "10110100"; x_in <= "01110101"; z_correct<="1101110101000100";
        when 13558 => y_in <= "10110100"; x_in <= "01110110"; z_correct<="1101110011111000";
        when 13559 => y_in <= "10110100"; x_in <= "01110111"; z_correct<="1101110010101100";
        when 13560 => y_in <= "10110100"; x_in <= "01111000"; z_correct<="1101110001100000";
        when 13561 => y_in <= "10110100"; x_in <= "01111001"; z_correct<="1101110000010100";
        when 13562 => y_in <= "10110100"; x_in <= "01111010"; z_correct<="1101101111001000";
        when 13563 => y_in <= "10110100"; x_in <= "01111011"; z_correct<="1101101101111100";
        when 13564 => y_in <= "10110100"; x_in <= "01111100"; z_correct<="1101101100110000";
        when 13565 => y_in <= "10110100"; x_in <= "01111101"; z_correct<="1101101011100100";
        when 13566 => y_in <= "10110100"; x_in <= "01111110"; z_correct<="1101101010011000";
        when 13567 => y_in <= "10110100"; x_in <= "01111111"; z_correct<="1101101001001100";
        when 13568 => y_in <= "10110101"; x_in <= "10000000"; z_correct<="0010010110000000";
        when 13569 => y_in <= "10110101"; x_in <= "10000001"; z_correct<="0010010100110101";
        when 13570 => y_in <= "10110101"; x_in <= "10000010"; z_correct<="0010010011101010";
        when 13571 => y_in <= "10110101"; x_in <= "10000011"; z_correct<="0010010010011111";
        when 13572 => y_in <= "10110101"; x_in <= "10000100"; z_correct<="0010010001010100";
        when 13573 => y_in <= "10110101"; x_in <= "10000101"; z_correct<="0010010000001001";
        when 13574 => y_in <= "10110101"; x_in <= "10000110"; z_correct<="0010001110111110";
        when 13575 => y_in <= "10110101"; x_in <= "10000111"; z_correct<="0010001101110011";
        when 13576 => y_in <= "10110101"; x_in <= "10001000"; z_correct<="0010001100101000";
        when 13577 => y_in <= "10110101"; x_in <= "10001001"; z_correct<="0010001011011101";
        when 13578 => y_in <= "10110101"; x_in <= "10001010"; z_correct<="0010001010010010";
        when 13579 => y_in <= "10110101"; x_in <= "10001011"; z_correct<="0010001001000111";
        when 13580 => y_in <= "10110101"; x_in <= "10001100"; z_correct<="0010000111111100";
        when 13581 => y_in <= "10110101"; x_in <= "10001101"; z_correct<="0010000110110001";
        when 13582 => y_in <= "10110101"; x_in <= "10001110"; z_correct<="0010000101100110";
        when 13583 => y_in <= "10110101"; x_in <= "10001111"; z_correct<="0010000100011011";
        when 13584 => y_in <= "10110101"; x_in <= "10010000"; z_correct<="0010000011010000";
        when 13585 => y_in <= "10110101"; x_in <= "10010001"; z_correct<="0010000010000101";
        when 13586 => y_in <= "10110101"; x_in <= "10010010"; z_correct<="0010000000111010";
        when 13587 => y_in <= "10110101"; x_in <= "10010011"; z_correct<="0001111111101111";
        when 13588 => y_in <= "10110101"; x_in <= "10010100"; z_correct<="0001111110100100";
        when 13589 => y_in <= "10110101"; x_in <= "10010101"; z_correct<="0001111101011001";
        when 13590 => y_in <= "10110101"; x_in <= "10010110"; z_correct<="0001111100001110";
        when 13591 => y_in <= "10110101"; x_in <= "10010111"; z_correct<="0001111011000011";
        when 13592 => y_in <= "10110101"; x_in <= "10011000"; z_correct<="0001111001111000";
        when 13593 => y_in <= "10110101"; x_in <= "10011001"; z_correct<="0001111000101101";
        when 13594 => y_in <= "10110101"; x_in <= "10011010"; z_correct<="0001110111100010";
        when 13595 => y_in <= "10110101"; x_in <= "10011011"; z_correct<="0001110110010111";
        when 13596 => y_in <= "10110101"; x_in <= "10011100"; z_correct<="0001110101001100";
        when 13597 => y_in <= "10110101"; x_in <= "10011101"; z_correct<="0001110100000001";
        when 13598 => y_in <= "10110101"; x_in <= "10011110"; z_correct<="0001110010110110";
        when 13599 => y_in <= "10110101"; x_in <= "10011111"; z_correct<="0001110001101011";
        when 13600 => y_in <= "10110101"; x_in <= "10100000"; z_correct<="0001110000100000";
        when 13601 => y_in <= "10110101"; x_in <= "10100001"; z_correct<="0001101111010101";
        when 13602 => y_in <= "10110101"; x_in <= "10100010"; z_correct<="0001101110001010";
        when 13603 => y_in <= "10110101"; x_in <= "10100011"; z_correct<="0001101100111111";
        when 13604 => y_in <= "10110101"; x_in <= "10100100"; z_correct<="0001101011110100";
        when 13605 => y_in <= "10110101"; x_in <= "10100101"; z_correct<="0001101010101001";
        when 13606 => y_in <= "10110101"; x_in <= "10100110"; z_correct<="0001101001011110";
        when 13607 => y_in <= "10110101"; x_in <= "10100111"; z_correct<="0001101000010011";
        when 13608 => y_in <= "10110101"; x_in <= "10101000"; z_correct<="0001100111001000";
        when 13609 => y_in <= "10110101"; x_in <= "10101001"; z_correct<="0001100101111101";
        when 13610 => y_in <= "10110101"; x_in <= "10101010"; z_correct<="0001100100110010";
        when 13611 => y_in <= "10110101"; x_in <= "10101011"; z_correct<="0001100011100111";
        when 13612 => y_in <= "10110101"; x_in <= "10101100"; z_correct<="0001100010011100";
        when 13613 => y_in <= "10110101"; x_in <= "10101101"; z_correct<="0001100001010001";
        when 13614 => y_in <= "10110101"; x_in <= "10101110"; z_correct<="0001100000000110";
        when 13615 => y_in <= "10110101"; x_in <= "10101111"; z_correct<="0001011110111011";
        when 13616 => y_in <= "10110101"; x_in <= "10110000"; z_correct<="0001011101110000";
        when 13617 => y_in <= "10110101"; x_in <= "10110001"; z_correct<="0001011100100101";
        when 13618 => y_in <= "10110101"; x_in <= "10110010"; z_correct<="0001011011011010";
        when 13619 => y_in <= "10110101"; x_in <= "10110011"; z_correct<="0001011010001111";
        when 13620 => y_in <= "10110101"; x_in <= "10110100"; z_correct<="0001011001000100";
        when 13621 => y_in <= "10110101"; x_in <= "10110101"; z_correct<="0001010111111001";
        when 13622 => y_in <= "10110101"; x_in <= "10110110"; z_correct<="0001010110101110";
        when 13623 => y_in <= "10110101"; x_in <= "10110111"; z_correct<="0001010101100011";
        when 13624 => y_in <= "10110101"; x_in <= "10111000"; z_correct<="0001010100011000";
        when 13625 => y_in <= "10110101"; x_in <= "10111001"; z_correct<="0001010011001101";
        when 13626 => y_in <= "10110101"; x_in <= "10111010"; z_correct<="0001010010000010";
        when 13627 => y_in <= "10110101"; x_in <= "10111011"; z_correct<="0001010000110111";
        when 13628 => y_in <= "10110101"; x_in <= "10111100"; z_correct<="0001001111101100";
        when 13629 => y_in <= "10110101"; x_in <= "10111101"; z_correct<="0001001110100001";
        when 13630 => y_in <= "10110101"; x_in <= "10111110"; z_correct<="0001001101010110";
        when 13631 => y_in <= "10110101"; x_in <= "10111111"; z_correct<="0001001100001011";
        when 13632 => y_in <= "10110101"; x_in <= "11000000"; z_correct<="0001001011000000";
        when 13633 => y_in <= "10110101"; x_in <= "11000001"; z_correct<="0001001001110101";
        when 13634 => y_in <= "10110101"; x_in <= "11000010"; z_correct<="0001001000101010";
        when 13635 => y_in <= "10110101"; x_in <= "11000011"; z_correct<="0001000111011111";
        when 13636 => y_in <= "10110101"; x_in <= "11000100"; z_correct<="0001000110010100";
        when 13637 => y_in <= "10110101"; x_in <= "11000101"; z_correct<="0001000101001001";
        when 13638 => y_in <= "10110101"; x_in <= "11000110"; z_correct<="0001000011111110";
        when 13639 => y_in <= "10110101"; x_in <= "11000111"; z_correct<="0001000010110011";
        when 13640 => y_in <= "10110101"; x_in <= "11001000"; z_correct<="0001000001101000";
        when 13641 => y_in <= "10110101"; x_in <= "11001001"; z_correct<="0001000000011101";
        when 13642 => y_in <= "10110101"; x_in <= "11001010"; z_correct<="0000111111010010";
        when 13643 => y_in <= "10110101"; x_in <= "11001011"; z_correct<="0000111110000111";
        when 13644 => y_in <= "10110101"; x_in <= "11001100"; z_correct<="0000111100111100";
        when 13645 => y_in <= "10110101"; x_in <= "11001101"; z_correct<="0000111011110001";
        when 13646 => y_in <= "10110101"; x_in <= "11001110"; z_correct<="0000111010100110";
        when 13647 => y_in <= "10110101"; x_in <= "11001111"; z_correct<="0000111001011011";
        when 13648 => y_in <= "10110101"; x_in <= "11010000"; z_correct<="0000111000010000";
        when 13649 => y_in <= "10110101"; x_in <= "11010001"; z_correct<="0000110111000101";
        when 13650 => y_in <= "10110101"; x_in <= "11010010"; z_correct<="0000110101111010";
        when 13651 => y_in <= "10110101"; x_in <= "11010011"; z_correct<="0000110100101111";
        when 13652 => y_in <= "10110101"; x_in <= "11010100"; z_correct<="0000110011100100";
        when 13653 => y_in <= "10110101"; x_in <= "11010101"; z_correct<="0000110010011001";
        when 13654 => y_in <= "10110101"; x_in <= "11010110"; z_correct<="0000110001001110";
        when 13655 => y_in <= "10110101"; x_in <= "11010111"; z_correct<="0000110000000011";
        when 13656 => y_in <= "10110101"; x_in <= "11011000"; z_correct<="0000101110111000";
        when 13657 => y_in <= "10110101"; x_in <= "11011001"; z_correct<="0000101101101101";
        when 13658 => y_in <= "10110101"; x_in <= "11011010"; z_correct<="0000101100100010";
        when 13659 => y_in <= "10110101"; x_in <= "11011011"; z_correct<="0000101011010111";
        when 13660 => y_in <= "10110101"; x_in <= "11011100"; z_correct<="0000101010001100";
        when 13661 => y_in <= "10110101"; x_in <= "11011101"; z_correct<="0000101001000001";
        when 13662 => y_in <= "10110101"; x_in <= "11011110"; z_correct<="0000100111110110";
        when 13663 => y_in <= "10110101"; x_in <= "11011111"; z_correct<="0000100110101011";
        when 13664 => y_in <= "10110101"; x_in <= "11100000"; z_correct<="0000100101100000";
        when 13665 => y_in <= "10110101"; x_in <= "11100001"; z_correct<="0000100100010101";
        when 13666 => y_in <= "10110101"; x_in <= "11100010"; z_correct<="0000100011001010";
        when 13667 => y_in <= "10110101"; x_in <= "11100011"; z_correct<="0000100001111111";
        when 13668 => y_in <= "10110101"; x_in <= "11100100"; z_correct<="0000100000110100";
        when 13669 => y_in <= "10110101"; x_in <= "11100101"; z_correct<="0000011111101001";
        when 13670 => y_in <= "10110101"; x_in <= "11100110"; z_correct<="0000011110011110";
        when 13671 => y_in <= "10110101"; x_in <= "11100111"; z_correct<="0000011101010011";
        when 13672 => y_in <= "10110101"; x_in <= "11101000"; z_correct<="0000011100001000";
        when 13673 => y_in <= "10110101"; x_in <= "11101001"; z_correct<="0000011010111101";
        when 13674 => y_in <= "10110101"; x_in <= "11101010"; z_correct<="0000011001110010";
        when 13675 => y_in <= "10110101"; x_in <= "11101011"; z_correct<="0000011000100111";
        when 13676 => y_in <= "10110101"; x_in <= "11101100"; z_correct<="0000010111011100";
        when 13677 => y_in <= "10110101"; x_in <= "11101101"; z_correct<="0000010110010001";
        when 13678 => y_in <= "10110101"; x_in <= "11101110"; z_correct<="0000010101000110";
        when 13679 => y_in <= "10110101"; x_in <= "11101111"; z_correct<="0000010011111011";
        when 13680 => y_in <= "10110101"; x_in <= "11110000"; z_correct<="0000010010110000";
        when 13681 => y_in <= "10110101"; x_in <= "11110001"; z_correct<="0000010001100101";
        when 13682 => y_in <= "10110101"; x_in <= "11110010"; z_correct<="0000010000011010";
        when 13683 => y_in <= "10110101"; x_in <= "11110011"; z_correct<="0000001111001111";
        when 13684 => y_in <= "10110101"; x_in <= "11110100"; z_correct<="0000001110000100";
        when 13685 => y_in <= "10110101"; x_in <= "11110101"; z_correct<="0000001100111001";
        when 13686 => y_in <= "10110101"; x_in <= "11110110"; z_correct<="0000001011101110";
        when 13687 => y_in <= "10110101"; x_in <= "11110111"; z_correct<="0000001010100011";
        when 13688 => y_in <= "10110101"; x_in <= "11111000"; z_correct<="0000001001011000";
        when 13689 => y_in <= "10110101"; x_in <= "11111001"; z_correct<="0000001000001101";
        when 13690 => y_in <= "10110101"; x_in <= "11111010"; z_correct<="0000000111000010";
        when 13691 => y_in <= "10110101"; x_in <= "11111011"; z_correct<="0000000101110111";
        when 13692 => y_in <= "10110101"; x_in <= "11111100"; z_correct<="0000000100101100";
        when 13693 => y_in <= "10110101"; x_in <= "11111101"; z_correct<="0000000011100001";
        when 13694 => y_in <= "10110101"; x_in <= "11111110"; z_correct<="0000000010010110";
        when 13695 => y_in <= "10110101"; x_in <= "11111111"; z_correct<="0000000001001011";
        when 13696 => y_in <= "10110101"; x_in <= "00000000"; z_correct<="0000000000000000";
        when 13697 => y_in <= "10110101"; x_in <= "00000001"; z_correct<="1111111110110101";
        when 13698 => y_in <= "10110101"; x_in <= "00000010"; z_correct<="1111111101101010";
        when 13699 => y_in <= "10110101"; x_in <= "00000011"; z_correct<="1111111100011111";
        when 13700 => y_in <= "10110101"; x_in <= "00000100"; z_correct<="1111111011010100";
        when 13701 => y_in <= "10110101"; x_in <= "00000101"; z_correct<="1111111010001001";
        when 13702 => y_in <= "10110101"; x_in <= "00000110"; z_correct<="1111111000111110";
        when 13703 => y_in <= "10110101"; x_in <= "00000111"; z_correct<="1111110111110011";
        when 13704 => y_in <= "10110101"; x_in <= "00001000"; z_correct<="1111110110101000";
        when 13705 => y_in <= "10110101"; x_in <= "00001001"; z_correct<="1111110101011101";
        when 13706 => y_in <= "10110101"; x_in <= "00001010"; z_correct<="1111110100010010";
        when 13707 => y_in <= "10110101"; x_in <= "00001011"; z_correct<="1111110011000111";
        when 13708 => y_in <= "10110101"; x_in <= "00001100"; z_correct<="1111110001111100";
        when 13709 => y_in <= "10110101"; x_in <= "00001101"; z_correct<="1111110000110001";
        when 13710 => y_in <= "10110101"; x_in <= "00001110"; z_correct<="1111101111100110";
        when 13711 => y_in <= "10110101"; x_in <= "00001111"; z_correct<="1111101110011011";
        when 13712 => y_in <= "10110101"; x_in <= "00010000"; z_correct<="1111101101010000";
        when 13713 => y_in <= "10110101"; x_in <= "00010001"; z_correct<="1111101100000101";
        when 13714 => y_in <= "10110101"; x_in <= "00010010"; z_correct<="1111101010111010";
        when 13715 => y_in <= "10110101"; x_in <= "00010011"; z_correct<="1111101001101111";
        when 13716 => y_in <= "10110101"; x_in <= "00010100"; z_correct<="1111101000100100";
        when 13717 => y_in <= "10110101"; x_in <= "00010101"; z_correct<="1111100111011001";
        when 13718 => y_in <= "10110101"; x_in <= "00010110"; z_correct<="1111100110001110";
        when 13719 => y_in <= "10110101"; x_in <= "00010111"; z_correct<="1111100101000011";
        when 13720 => y_in <= "10110101"; x_in <= "00011000"; z_correct<="1111100011111000";
        when 13721 => y_in <= "10110101"; x_in <= "00011001"; z_correct<="1111100010101101";
        when 13722 => y_in <= "10110101"; x_in <= "00011010"; z_correct<="1111100001100010";
        when 13723 => y_in <= "10110101"; x_in <= "00011011"; z_correct<="1111100000010111";
        when 13724 => y_in <= "10110101"; x_in <= "00011100"; z_correct<="1111011111001100";
        when 13725 => y_in <= "10110101"; x_in <= "00011101"; z_correct<="1111011110000001";
        when 13726 => y_in <= "10110101"; x_in <= "00011110"; z_correct<="1111011100110110";
        when 13727 => y_in <= "10110101"; x_in <= "00011111"; z_correct<="1111011011101011";
        when 13728 => y_in <= "10110101"; x_in <= "00100000"; z_correct<="1111011010100000";
        when 13729 => y_in <= "10110101"; x_in <= "00100001"; z_correct<="1111011001010101";
        when 13730 => y_in <= "10110101"; x_in <= "00100010"; z_correct<="1111011000001010";
        when 13731 => y_in <= "10110101"; x_in <= "00100011"; z_correct<="1111010110111111";
        when 13732 => y_in <= "10110101"; x_in <= "00100100"; z_correct<="1111010101110100";
        when 13733 => y_in <= "10110101"; x_in <= "00100101"; z_correct<="1111010100101001";
        when 13734 => y_in <= "10110101"; x_in <= "00100110"; z_correct<="1111010011011110";
        when 13735 => y_in <= "10110101"; x_in <= "00100111"; z_correct<="1111010010010011";
        when 13736 => y_in <= "10110101"; x_in <= "00101000"; z_correct<="1111010001001000";
        when 13737 => y_in <= "10110101"; x_in <= "00101001"; z_correct<="1111001111111101";
        when 13738 => y_in <= "10110101"; x_in <= "00101010"; z_correct<="1111001110110010";
        when 13739 => y_in <= "10110101"; x_in <= "00101011"; z_correct<="1111001101100111";
        when 13740 => y_in <= "10110101"; x_in <= "00101100"; z_correct<="1111001100011100";
        when 13741 => y_in <= "10110101"; x_in <= "00101101"; z_correct<="1111001011010001";
        when 13742 => y_in <= "10110101"; x_in <= "00101110"; z_correct<="1111001010000110";
        when 13743 => y_in <= "10110101"; x_in <= "00101111"; z_correct<="1111001000111011";
        when 13744 => y_in <= "10110101"; x_in <= "00110000"; z_correct<="1111000111110000";
        when 13745 => y_in <= "10110101"; x_in <= "00110001"; z_correct<="1111000110100101";
        when 13746 => y_in <= "10110101"; x_in <= "00110010"; z_correct<="1111000101011010";
        when 13747 => y_in <= "10110101"; x_in <= "00110011"; z_correct<="1111000100001111";
        when 13748 => y_in <= "10110101"; x_in <= "00110100"; z_correct<="1111000011000100";
        when 13749 => y_in <= "10110101"; x_in <= "00110101"; z_correct<="1111000001111001";
        when 13750 => y_in <= "10110101"; x_in <= "00110110"; z_correct<="1111000000101110";
        when 13751 => y_in <= "10110101"; x_in <= "00110111"; z_correct<="1110111111100011";
        when 13752 => y_in <= "10110101"; x_in <= "00111000"; z_correct<="1110111110011000";
        when 13753 => y_in <= "10110101"; x_in <= "00111001"; z_correct<="1110111101001101";
        when 13754 => y_in <= "10110101"; x_in <= "00111010"; z_correct<="1110111100000010";
        when 13755 => y_in <= "10110101"; x_in <= "00111011"; z_correct<="1110111010110111";
        when 13756 => y_in <= "10110101"; x_in <= "00111100"; z_correct<="1110111001101100";
        when 13757 => y_in <= "10110101"; x_in <= "00111101"; z_correct<="1110111000100001";
        when 13758 => y_in <= "10110101"; x_in <= "00111110"; z_correct<="1110110111010110";
        when 13759 => y_in <= "10110101"; x_in <= "00111111"; z_correct<="1110110110001011";
        when 13760 => y_in <= "10110101"; x_in <= "01000000"; z_correct<="1110110101000000";
        when 13761 => y_in <= "10110101"; x_in <= "01000001"; z_correct<="1110110011110101";
        when 13762 => y_in <= "10110101"; x_in <= "01000010"; z_correct<="1110110010101010";
        when 13763 => y_in <= "10110101"; x_in <= "01000011"; z_correct<="1110110001011111";
        when 13764 => y_in <= "10110101"; x_in <= "01000100"; z_correct<="1110110000010100";
        when 13765 => y_in <= "10110101"; x_in <= "01000101"; z_correct<="1110101111001001";
        when 13766 => y_in <= "10110101"; x_in <= "01000110"; z_correct<="1110101101111110";
        when 13767 => y_in <= "10110101"; x_in <= "01000111"; z_correct<="1110101100110011";
        when 13768 => y_in <= "10110101"; x_in <= "01001000"; z_correct<="1110101011101000";
        when 13769 => y_in <= "10110101"; x_in <= "01001001"; z_correct<="1110101010011101";
        when 13770 => y_in <= "10110101"; x_in <= "01001010"; z_correct<="1110101001010010";
        when 13771 => y_in <= "10110101"; x_in <= "01001011"; z_correct<="1110101000000111";
        when 13772 => y_in <= "10110101"; x_in <= "01001100"; z_correct<="1110100110111100";
        when 13773 => y_in <= "10110101"; x_in <= "01001101"; z_correct<="1110100101110001";
        when 13774 => y_in <= "10110101"; x_in <= "01001110"; z_correct<="1110100100100110";
        when 13775 => y_in <= "10110101"; x_in <= "01001111"; z_correct<="1110100011011011";
        when 13776 => y_in <= "10110101"; x_in <= "01010000"; z_correct<="1110100010010000";
        when 13777 => y_in <= "10110101"; x_in <= "01010001"; z_correct<="1110100001000101";
        when 13778 => y_in <= "10110101"; x_in <= "01010010"; z_correct<="1110011111111010";
        when 13779 => y_in <= "10110101"; x_in <= "01010011"; z_correct<="1110011110101111";
        when 13780 => y_in <= "10110101"; x_in <= "01010100"; z_correct<="1110011101100100";
        when 13781 => y_in <= "10110101"; x_in <= "01010101"; z_correct<="1110011100011001";
        when 13782 => y_in <= "10110101"; x_in <= "01010110"; z_correct<="1110011011001110";
        when 13783 => y_in <= "10110101"; x_in <= "01010111"; z_correct<="1110011010000011";
        when 13784 => y_in <= "10110101"; x_in <= "01011000"; z_correct<="1110011000111000";
        when 13785 => y_in <= "10110101"; x_in <= "01011001"; z_correct<="1110010111101101";
        when 13786 => y_in <= "10110101"; x_in <= "01011010"; z_correct<="1110010110100010";
        when 13787 => y_in <= "10110101"; x_in <= "01011011"; z_correct<="1110010101010111";
        when 13788 => y_in <= "10110101"; x_in <= "01011100"; z_correct<="1110010100001100";
        when 13789 => y_in <= "10110101"; x_in <= "01011101"; z_correct<="1110010011000001";
        when 13790 => y_in <= "10110101"; x_in <= "01011110"; z_correct<="1110010001110110";
        when 13791 => y_in <= "10110101"; x_in <= "01011111"; z_correct<="1110010000101011";
        when 13792 => y_in <= "10110101"; x_in <= "01100000"; z_correct<="1110001111100000";
        when 13793 => y_in <= "10110101"; x_in <= "01100001"; z_correct<="1110001110010101";
        when 13794 => y_in <= "10110101"; x_in <= "01100010"; z_correct<="1110001101001010";
        when 13795 => y_in <= "10110101"; x_in <= "01100011"; z_correct<="1110001011111111";
        when 13796 => y_in <= "10110101"; x_in <= "01100100"; z_correct<="1110001010110100";
        when 13797 => y_in <= "10110101"; x_in <= "01100101"; z_correct<="1110001001101001";
        when 13798 => y_in <= "10110101"; x_in <= "01100110"; z_correct<="1110001000011110";
        when 13799 => y_in <= "10110101"; x_in <= "01100111"; z_correct<="1110000111010011";
        when 13800 => y_in <= "10110101"; x_in <= "01101000"; z_correct<="1110000110001000";
        when 13801 => y_in <= "10110101"; x_in <= "01101001"; z_correct<="1110000100111101";
        when 13802 => y_in <= "10110101"; x_in <= "01101010"; z_correct<="1110000011110010";
        when 13803 => y_in <= "10110101"; x_in <= "01101011"; z_correct<="1110000010100111";
        when 13804 => y_in <= "10110101"; x_in <= "01101100"; z_correct<="1110000001011100";
        when 13805 => y_in <= "10110101"; x_in <= "01101101"; z_correct<="1110000000010001";
        when 13806 => y_in <= "10110101"; x_in <= "01101110"; z_correct<="1101111111000110";
        when 13807 => y_in <= "10110101"; x_in <= "01101111"; z_correct<="1101111101111011";
        when 13808 => y_in <= "10110101"; x_in <= "01110000"; z_correct<="1101111100110000";
        when 13809 => y_in <= "10110101"; x_in <= "01110001"; z_correct<="1101111011100101";
        when 13810 => y_in <= "10110101"; x_in <= "01110010"; z_correct<="1101111010011010";
        when 13811 => y_in <= "10110101"; x_in <= "01110011"; z_correct<="1101111001001111";
        when 13812 => y_in <= "10110101"; x_in <= "01110100"; z_correct<="1101111000000100";
        when 13813 => y_in <= "10110101"; x_in <= "01110101"; z_correct<="1101110110111001";
        when 13814 => y_in <= "10110101"; x_in <= "01110110"; z_correct<="1101110101101110";
        when 13815 => y_in <= "10110101"; x_in <= "01110111"; z_correct<="1101110100100011";
        when 13816 => y_in <= "10110101"; x_in <= "01111000"; z_correct<="1101110011011000";
        when 13817 => y_in <= "10110101"; x_in <= "01111001"; z_correct<="1101110010001101";
        when 13818 => y_in <= "10110101"; x_in <= "01111010"; z_correct<="1101110001000010";
        when 13819 => y_in <= "10110101"; x_in <= "01111011"; z_correct<="1101101111110111";
        when 13820 => y_in <= "10110101"; x_in <= "01111100"; z_correct<="1101101110101100";
        when 13821 => y_in <= "10110101"; x_in <= "01111101"; z_correct<="1101101101100001";
        when 13822 => y_in <= "10110101"; x_in <= "01111110"; z_correct<="1101101100010110";
        when 13823 => y_in <= "10110101"; x_in <= "01111111"; z_correct<="1101101011001011";
        when 13824 => y_in <= "10110110"; x_in <= "10000000"; z_correct<="0010010100000000";
        when 13825 => y_in <= "10110110"; x_in <= "10000001"; z_correct<="0010010010110110";
        when 13826 => y_in <= "10110110"; x_in <= "10000010"; z_correct<="0010010001101100";
        when 13827 => y_in <= "10110110"; x_in <= "10000011"; z_correct<="0010010000100010";
        when 13828 => y_in <= "10110110"; x_in <= "10000100"; z_correct<="0010001111011000";
        when 13829 => y_in <= "10110110"; x_in <= "10000101"; z_correct<="0010001110001110";
        when 13830 => y_in <= "10110110"; x_in <= "10000110"; z_correct<="0010001101000100";
        when 13831 => y_in <= "10110110"; x_in <= "10000111"; z_correct<="0010001011111010";
        when 13832 => y_in <= "10110110"; x_in <= "10001000"; z_correct<="0010001010110000";
        when 13833 => y_in <= "10110110"; x_in <= "10001001"; z_correct<="0010001001100110";
        when 13834 => y_in <= "10110110"; x_in <= "10001010"; z_correct<="0010001000011100";
        when 13835 => y_in <= "10110110"; x_in <= "10001011"; z_correct<="0010000111010010";
        when 13836 => y_in <= "10110110"; x_in <= "10001100"; z_correct<="0010000110001000";
        when 13837 => y_in <= "10110110"; x_in <= "10001101"; z_correct<="0010000100111110";
        when 13838 => y_in <= "10110110"; x_in <= "10001110"; z_correct<="0010000011110100";
        when 13839 => y_in <= "10110110"; x_in <= "10001111"; z_correct<="0010000010101010";
        when 13840 => y_in <= "10110110"; x_in <= "10010000"; z_correct<="0010000001100000";
        when 13841 => y_in <= "10110110"; x_in <= "10010001"; z_correct<="0010000000010110";
        when 13842 => y_in <= "10110110"; x_in <= "10010010"; z_correct<="0001111111001100";
        when 13843 => y_in <= "10110110"; x_in <= "10010011"; z_correct<="0001111110000010";
        when 13844 => y_in <= "10110110"; x_in <= "10010100"; z_correct<="0001111100111000";
        when 13845 => y_in <= "10110110"; x_in <= "10010101"; z_correct<="0001111011101110";
        when 13846 => y_in <= "10110110"; x_in <= "10010110"; z_correct<="0001111010100100";
        when 13847 => y_in <= "10110110"; x_in <= "10010111"; z_correct<="0001111001011010";
        when 13848 => y_in <= "10110110"; x_in <= "10011000"; z_correct<="0001111000010000";
        when 13849 => y_in <= "10110110"; x_in <= "10011001"; z_correct<="0001110111000110";
        when 13850 => y_in <= "10110110"; x_in <= "10011010"; z_correct<="0001110101111100";
        when 13851 => y_in <= "10110110"; x_in <= "10011011"; z_correct<="0001110100110010";
        when 13852 => y_in <= "10110110"; x_in <= "10011100"; z_correct<="0001110011101000";
        when 13853 => y_in <= "10110110"; x_in <= "10011101"; z_correct<="0001110010011110";
        when 13854 => y_in <= "10110110"; x_in <= "10011110"; z_correct<="0001110001010100";
        when 13855 => y_in <= "10110110"; x_in <= "10011111"; z_correct<="0001110000001010";
        when 13856 => y_in <= "10110110"; x_in <= "10100000"; z_correct<="0001101111000000";
        when 13857 => y_in <= "10110110"; x_in <= "10100001"; z_correct<="0001101101110110";
        when 13858 => y_in <= "10110110"; x_in <= "10100010"; z_correct<="0001101100101100";
        when 13859 => y_in <= "10110110"; x_in <= "10100011"; z_correct<="0001101011100010";
        when 13860 => y_in <= "10110110"; x_in <= "10100100"; z_correct<="0001101010011000";
        when 13861 => y_in <= "10110110"; x_in <= "10100101"; z_correct<="0001101001001110";
        when 13862 => y_in <= "10110110"; x_in <= "10100110"; z_correct<="0001101000000100";
        when 13863 => y_in <= "10110110"; x_in <= "10100111"; z_correct<="0001100110111010";
        when 13864 => y_in <= "10110110"; x_in <= "10101000"; z_correct<="0001100101110000";
        when 13865 => y_in <= "10110110"; x_in <= "10101001"; z_correct<="0001100100100110";
        when 13866 => y_in <= "10110110"; x_in <= "10101010"; z_correct<="0001100011011100";
        when 13867 => y_in <= "10110110"; x_in <= "10101011"; z_correct<="0001100010010010";
        when 13868 => y_in <= "10110110"; x_in <= "10101100"; z_correct<="0001100001001000";
        when 13869 => y_in <= "10110110"; x_in <= "10101101"; z_correct<="0001011111111110";
        when 13870 => y_in <= "10110110"; x_in <= "10101110"; z_correct<="0001011110110100";
        when 13871 => y_in <= "10110110"; x_in <= "10101111"; z_correct<="0001011101101010";
        when 13872 => y_in <= "10110110"; x_in <= "10110000"; z_correct<="0001011100100000";
        when 13873 => y_in <= "10110110"; x_in <= "10110001"; z_correct<="0001011011010110";
        when 13874 => y_in <= "10110110"; x_in <= "10110010"; z_correct<="0001011010001100";
        when 13875 => y_in <= "10110110"; x_in <= "10110011"; z_correct<="0001011001000010";
        when 13876 => y_in <= "10110110"; x_in <= "10110100"; z_correct<="0001010111111000";
        when 13877 => y_in <= "10110110"; x_in <= "10110101"; z_correct<="0001010110101110";
        when 13878 => y_in <= "10110110"; x_in <= "10110110"; z_correct<="0001010101100100";
        when 13879 => y_in <= "10110110"; x_in <= "10110111"; z_correct<="0001010100011010";
        when 13880 => y_in <= "10110110"; x_in <= "10111000"; z_correct<="0001010011010000";
        when 13881 => y_in <= "10110110"; x_in <= "10111001"; z_correct<="0001010010000110";
        when 13882 => y_in <= "10110110"; x_in <= "10111010"; z_correct<="0001010000111100";
        when 13883 => y_in <= "10110110"; x_in <= "10111011"; z_correct<="0001001111110010";
        when 13884 => y_in <= "10110110"; x_in <= "10111100"; z_correct<="0001001110101000";
        when 13885 => y_in <= "10110110"; x_in <= "10111101"; z_correct<="0001001101011110";
        when 13886 => y_in <= "10110110"; x_in <= "10111110"; z_correct<="0001001100010100";
        when 13887 => y_in <= "10110110"; x_in <= "10111111"; z_correct<="0001001011001010";
        when 13888 => y_in <= "10110110"; x_in <= "11000000"; z_correct<="0001001010000000";
        when 13889 => y_in <= "10110110"; x_in <= "11000001"; z_correct<="0001001000110110";

        when (13895) =>   Testing <= False;
        when others => null;
     end case;
	 if (z_out = z_correct) then diff <= '0'; else diff <= '1'; end if;
     count:= count + 1;
   end process Test_Proc;
end booth2_tbn8;
