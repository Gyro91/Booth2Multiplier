							  

library IEEE;
use IEEE.std_logic_1164.all;

entity booth2_tbnm is

end booth2_tbnm;

-- Test Booth Multiplier with N!=M

architecture booth2_tbnm of booth2_tbnm is
	component Booth2Multiplier
  	generic(N : integer := 4; 
            M : integer := 4   
       );
	port (
	x : in  std_logic_vector(N-1 downto 0); 	-- x is the multiplicand
	y : in  std_logic_vector(M-1 downto 0);		-- y is the multiplier
	z : out	std_logic_vector(N+M-1 downto 0)	-- z is the result of the multiplication
		);
	end component; 
	
   constant MckPer  :  time     := 200 ns;  
	   
   signal   clk  : std_logic := '0';
   signal   x_in   	: std_logic_VECTOR (5 downto 0):="000000";
   signal   y_in    : std_logic_VECTOR (3 downto 0):="0000";	
   signal   z_out   : std_logic_VECTOR (9 downto 0):="0000000000";
   signal clk_cycle : integer;
   signal Testing: boolean := True;	
   signal z_correct   : std_logic_VECTOR (9 downto 0):="0000000000";
   signal 	diff		: std_logic := '0';
begin 			 
	I: Booth2Multiplier generic map(N=>6, M=>4)
		port map(x=>x_in,y=>y_in, z=>z_out);
				
		clk <= not clk after MckPer/2 when Testing else '0';

   Test_Proc: process(clk)
   variable count: INTEGER:= 0;
   
   begin
     clk_cycle <= (count+1)/2;

     case clk_cycle is

        when 0 => y_in <= "1000"; x_in <= "100000"; z_correct<="0100000000";
        when 1 => y_in <= "1001"; x_in <= "100000"; z_correct<="0011100000";
        when 2 => y_in <= "1010"; x_in <= "100000"; z_correct<="0011000000";
        when 3 => y_in <= "1011"; x_in <= "100000"; z_correct<="0010100000";
        when 4 => y_in <= "1100"; x_in <= "100000"; z_correct<="0010000000";
        when 5 => y_in <= "1101"; x_in <= "100000"; z_correct<="0001100000";
        when 6 => y_in <= "1110"; x_in <= "100000"; z_correct<="0001000000";
        when 7 => y_in <= "1111"; x_in <= "100000"; z_correct<="0000100000";
        when 8 => y_in <= "0000"; x_in <= "100000"; z_correct<="0000000000";
        when 9 => y_in <= "0001"; x_in <= "100000"; z_correct<="1111100000";
        when 10 => y_in <= "0010"; x_in <= "100000"; z_correct<="1111000000";
        when 11 => y_in <= "0011"; x_in <= "100000"; z_correct<="1110100000";
        when 12 => y_in <= "0100"; x_in <= "100000"; z_correct<="1110000000";
        when 13 => y_in <= "0101"; x_in <= "100000"; z_correct<="1101100000";
        when 14 => y_in <= "0110"; x_in <= "100000"; z_correct<="1101000000";
        when 15 => y_in <= "0111"; x_in <= "100000"; z_correct<="1100100000";
        when 16 => y_in <= "1000"; x_in <= "100001"; z_correct<="0011111000";
        when 17 => y_in <= "1001"; x_in <= "100001"; z_correct<="0011011001";
        when 18 => y_in <= "1010"; x_in <= "100001"; z_correct<="0010111010";
        when 19 => y_in <= "1011"; x_in <= "100001"; z_correct<="0010011011";
        when 20 => y_in <= "1100"; x_in <= "100001"; z_correct<="0001111100";
        when 21 => y_in <= "1101"; x_in <= "100001"; z_correct<="0001011101";
        when 22 => y_in <= "1110"; x_in <= "100001"; z_correct<="0000111110";
        when 23 => y_in <= "1111"; x_in <= "100001"; z_correct<="0000011111";
        when 24 => y_in <= "0000"; x_in <= "100001"; z_correct<="0000000000";
        when 25 => y_in <= "0001"; x_in <= "100001"; z_correct<="1111100001";
        when 26 => y_in <= "0010"; x_in <= "100001"; z_correct<="1111000010";
        when 27 => y_in <= "0011"; x_in <= "100001"; z_correct<="1110100011";
        when 28 => y_in <= "0100"; x_in <= "100001"; z_correct<="1110000100";
        when 29 => y_in <= "0101"; x_in <= "100001"; z_correct<="1101100101";
        when 30 => y_in <= "0110"; x_in <= "100001"; z_correct<="1101000110";
        when 31 => y_in <= "0111"; x_in <= "100001"; z_correct<="1100100111";
        when 32 => y_in <= "1000"; x_in <= "100010"; z_correct<="0011110000";
        when 33 => y_in <= "1001"; x_in <= "100010"; z_correct<="0011010010";
        when 34 => y_in <= "1010"; x_in <= "100010"; z_correct<="0010110100";
        when 35 => y_in <= "1011"; x_in <= "100010"; z_correct<="0010010110";
        when 36 => y_in <= "1100"; x_in <= "100010"; z_correct<="0001111000";
        when 37 => y_in <= "1101"; x_in <= "100010"; z_correct<="0001011010";
        when 38 => y_in <= "1110"; x_in <= "100010"; z_correct<="0000111100";
        when 39 => y_in <= "1111"; x_in <= "100010"; z_correct<="0000011110";
        when 40 => y_in <= "0000"; x_in <= "100010"; z_correct<="0000000000";
        when 41 => y_in <= "0001"; x_in <= "100010"; z_correct<="1111100010";
        when 42 => y_in <= "0010"; x_in <= "100010"; z_correct<="1111000100";
        when 43 => y_in <= "0011"; x_in <= "100010"; z_correct<="1110100110";
        when 44 => y_in <= "0100"; x_in <= "100010"; z_correct<="1110001000";
        when 45 => y_in <= "0101"; x_in <= "100010"; z_correct<="1101101010";
        when 46 => y_in <= "0110"; x_in <= "100010"; z_correct<="1101001100";
        when 47 => y_in <= "0111"; x_in <= "100010"; z_correct<="1100101110";
        when 48 => y_in <= "1000"; x_in <= "100011"; z_correct<="0011101000";
        when 49 => y_in <= "1001"; x_in <= "100011"; z_correct<="0011001011";
        when 50 => y_in <= "1010"; x_in <= "100011"; z_correct<="0010101110";
        when 51 => y_in <= "1011"; x_in <= "100011"; z_correct<="0010010001";
        when 52 => y_in <= "1100"; x_in <= "100011"; z_correct<="0001110100";
        when 53 => y_in <= "1101"; x_in <= "100011"; z_correct<="0001010111";
        when 54 => y_in <= "1110"; x_in <= "100011"; z_correct<="0000111010";
        when 55 => y_in <= "1111"; x_in <= "100011"; z_correct<="0000011101";
        when 56 => y_in <= "0000"; x_in <= "100011"; z_correct<="0000000000";
        when 57 => y_in <= "0001"; x_in <= "100011"; z_correct<="1111100011";
        when 58 => y_in <= "0010"; x_in <= "100011"; z_correct<="1111000110";
        when 59 => y_in <= "0011"; x_in <= "100011"; z_correct<="1110101001";
        when 60 => y_in <= "0100"; x_in <= "100011"; z_correct<="1110001100";
        when 61 => y_in <= "0101"; x_in <= "100011"; z_correct<="1101101111";
        when 62 => y_in <= "0110"; x_in <= "100011"; z_correct<="1101010010";
        when 63 => y_in <= "0111"; x_in <= "100011"; z_correct<="1100110101";
        when 64 => y_in <= "1000"; x_in <= "100100"; z_correct<="0011100000";
        when 65 => y_in <= "1001"; x_in <= "100100"; z_correct<="0011000100";
        when 66 => y_in <= "1010"; x_in <= "100100"; z_correct<="0010101000";
        when 67 => y_in <= "1011"; x_in <= "100100"; z_correct<="0010001100";
        when 68 => y_in <= "1100"; x_in <= "100100"; z_correct<="0001110000";
        when 69 => y_in <= "1101"; x_in <= "100100"; z_correct<="0001010100";
        when 70 => y_in <= "1110"; x_in <= "100100"; z_correct<="0000111000";
        when 71 => y_in <= "1111"; x_in <= "100100"; z_correct<="0000011100";
        when 72 => y_in <= "0000"; x_in <= "100100"; z_correct<="0000000000";
        when 73 => y_in <= "0001"; x_in <= "100100"; z_correct<="1111100100";
        when 74 => y_in <= "0010"; x_in <= "100100"; z_correct<="1111001000";
        when 75 => y_in <= "0011"; x_in <= "100100"; z_correct<="1110101100";
        when 76 => y_in <= "0100"; x_in <= "100100"; z_correct<="1110010000";
        when 77 => y_in <= "0101"; x_in <= "100100"; z_correct<="1101110100";
        when 78 => y_in <= "0110"; x_in <= "100100"; z_correct<="1101011000";
        when 79 => y_in <= "0111"; x_in <= "100100"; z_correct<="1100111100";
        when 80 => y_in <= "1000"; x_in <= "100101"; z_correct<="0011011000";
        when 81 => y_in <= "1001"; x_in <= "100101"; z_correct<="0010111101";
        when 82 => y_in <= "1010"; x_in <= "100101"; z_correct<="0010100010";
        when 83 => y_in <= "1011"; x_in <= "100101"; z_correct<="0010000111";
        when 84 => y_in <= "1100"; x_in <= "100101"; z_correct<="0001101100";
        when 85 => y_in <= "1101"; x_in <= "100101"; z_correct<="0001010001";
        when 86 => y_in <= "1110"; x_in <= "100101"; z_correct<="0000110110";
        when 87 => y_in <= "1111"; x_in <= "100101"; z_correct<="0000011011";
        when 88 => y_in <= "0000"; x_in <= "100101"; z_correct<="0000000000";
        when 89 => y_in <= "0001"; x_in <= "100101"; z_correct<="1111100101";
        when 90 => y_in <= "0010"; x_in <= "100101"; z_correct<="1111001010";
        when 91 => y_in <= "0011"; x_in <= "100101"; z_correct<="1110101111";
        when 92 => y_in <= "0100"; x_in <= "100101"; z_correct<="1110010100";
        when 93 => y_in <= "0101"; x_in <= "100101"; z_correct<="1101111001";
        when 94 => y_in <= "0110"; x_in <= "100101"; z_correct<="1101011110";
        when 95 => y_in <= "0111"; x_in <= "100101"; z_correct<="1101000011";
        when 96 => y_in <= "1000"; x_in <= "100110"; z_correct<="0011010000";
        when 97 => y_in <= "1001"; x_in <= "100110"; z_correct<="0010110110";
        when 98 => y_in <= "1010"; x_in <= "100110"; z_correct<="0010011100";
        when 99 => y_in <= "1011"; x_in <= "100110"; z_correct<="0010000010";
        when 100 => y_in <= "1100"; x_in <= "100110"; z_correct<="0001101000";
        when 101 => y_in <= "1101"; x_in <= "100110"; z_correct<="0001001110";
        when 102 => y_in <= "1110"; x_in <= "100110"; z_correct<="0000110100";
        when 103 => y_in <= "1111"; x_in <= "100110"; z_correct<="0000011010";
        when 104 => y_in <= "0000"; x_in <= "100110"; z_correct<="0000000000";
        when 105 => y_in <= "0001"; x_in <= "100110"; z_correct<="1111100110";
        when 106 => y_in <= "0010"; x_in <= "100110"; z_correct<="1111001100";
        when 107 => y_in <= "0011"; x_in <= "100110"; z_correct<="1110110010";
        when 108 => y_in <= "0100"; x_in <= "100110"; z_correct<="1110011000";
        when 109 => y_in <= "0101"; x_in <= "100110"; z_correct<="1101111110";
        when 110 => y_in <= "0110"; x_in <= "100110"; z_correct<="1101100100";
        when 111 => y_in <= "0111"; x_in <= "100110"; z_correct<="1101001010";
        when 112 => y_in <= "1000"; x_in <= "100111"; z_correct<="0011001000";
        when 113 => y_in <= "1001"; x_in <= "100111"; z_correct<="0010101111";
        when 114 => y_in <= "1010"; x_in <= "100111"; z_correct<="0010010110";
        when 115 => y_in <= "1011"; x_in <= "100111"; z_correct<="0001111101";
        when 116 => y_in <= "1100"; x_in <= "100111"; z_correct<="0001100100";
        when 117 => y_in <= "1101"; x_in <= "100111"; z_correct<="0001001011";
        when 118 => y_in <= "1110"; x_in <= "100111"; z_correct<="0000110010";
        when 119 => y_in <= "1111"; x_in <= "100111"; z_correct<="0000011001";
        when 120 => y_in <= "0000"; x_in <= "100111"; z_correct<="0000000000";
        when 121 => y_in <= "0001"; x_in <= "100111"; z_correct<="1111100111";
        when 122 => y_in <= "0010"; x_in <= "100111"; z_correct<="1111001110";
        when 123 => y_in <= "0011"; x_in <= "100111"; z_correct<="1110110101";
        when 124 => y_in <= "0100"; x_in <= "100111"; z_correct<="1110011100";
        when 125 => y_in <= "0101"; x_in <= "100111"; z_correct<="1110000011";
        when 126 => y_in <= "0110"; x_in <= "100111"; z_correct<="1101101010";
        when 127 => y_in <= "0111"; x_in <= "100111"; z_correct<="1101010001";
        when 128 => y_in <= "1000"; x_in <= "101000"; z_correct<="0011000000";
        when 129 => y_in <= "1001"; x_in <= "101000"; z_correct<="0010101000";
        when 130 => y_in <= "1010"; x_in <= "101000"; z_correct<="0010010000";
        when 131 => y_in <= "1011"; x_in <= "101000"; z_correct<="0001111000";
        when 132 => y_in <= "1100"; x_in <= "101000"; z_correct<="0001100000";
        when 133 => y_in <= "1101"; x_in <= "101000"; z_correct<="0001001000";
        when 134 => y_in <= "1110"; x_in <= "101000"; z_correct<="0000110000";
        when 135 => y_in <= "1111"; x_in <= "101000"; z_correct<="0000011000";
        when 136 => y_in <= "0000"; x_in <= "101000"; z_correct<="0000000000";
        when 137 => y_in <= "0001"; x_in <= "101000"; z_correct<="1111101000";
        when 138 => y_in <= "0010"; x_in <= "101000"; z_correct<="1111010000";
        when 139 => y_in <= "0011"; x_in <= "101000"; z_correct<="1110111000";
        when 140 => y_in <= "0100"; x_in <= "101000"; z_correct<="1110100000";
        when 141 => y_in <= "0101"; x_in <= "101000"; z_correct<="1110001000";
        when 142 => y_in <= "0110"; x_in <= "101000"; z_correct<="1101110000";
        when 143 => y_in <= "0111"; x_in <= "101000"; z_correct<="1101011000";
        when 144 => y_in <= "1000"; x_in <= "101001"; z_correct<="0010111000";
        when 145 => y_in <= "1001"; x_in <= "101001"; z_correct<="0010100001";
        when 146 => y_in <= "1010"; x_in <= "101001"; z_correct<="0010001010";
        when 147 => y_in <= "1011"; x_in <= "101001"; z_correct<="0001110011";
        when 148 => y_in <= "1100"; x_in <= "101001"; z_correct<="0001011100";
        when 149 => y_in <= "1101"; x_in <= "101001"; z_correct<="0001000101";
        when 150 => y_in <= "1110"; x_in <= "101001"; z_correct<="0000101110";
        when 151 => y_in <= "1111"; x_in <= "101001"; z_correct<="0000010111";
        when 152 => y_in <= "0000"; x_in <= "101001"; z_correct<="0000000000";
        when 153 => y_in <= "0001"; x_in <= "101001"; z_correct<="1111101001";
        when 154 => y_in <= "0010"; x_in <= "101001"; z_correct<="1111010010";
        when 155 => y_in <= "0011"; x_in <= "101001"; z_correct<="1110111011";
        when 156 => y_in <= "0100"; x_in <= "101001"; z_correct<="1110100100";
        when 157 => y_in <= "0101"; x_in <= "101001"; z_correct<="1110001101";
        when 158 => y_in <= "0110"; x_in <= "101001"; z_correct<="1101110110";
        when 159 => y_in <= "0111"; x_in <= "101001"; z_correct<="1101011111";
        when 160 => y_in <= "1000"; x_in <= "101010"; z_correct<="0010110000";
        when 161 => y_in <= "1001"; x_in <= "101010"; z_correct<="0010011010";
        when 162 => y_in <= "1010"; x_in <= "101010"; z_correct<="0010000100";
        when 163 => y_in <= "1011"; x_in <= "101010"; z_correct<="0001101110";
        when 164 => y_in <= "1100"; x_in <= "101010"; z_correct<="0001011000";
        when 165 => y_in <= "1101"; x_in <= "101010"; z_correct<="0001000010";
        when 166 => y_in <= "1110"; x_in <= "101010"; z_correct<="0000101100";
        when 167 => y_in <= "1111"; x_in <= "101010"; z_correct<="0000010110";
        when 168 => y_in <= "0000"; x_in <= "101010"; z_correct<="0000000000";
        when 169 => y_in <= "0001"; x_in <= "101010"; z_correct<="1111101010";
        when 170 => y_in <= "0010"; x_in <= "101010"; z_correct<="1111010100";
        when 171 => y_in <= "0011"; x_in <= "101010"; z_correct<="1110111110";
        when 172 => y_in <= "0100"; x_in <= "101010"; z_correct<="1110101000";
        when 173 => y_in <= "0101"; x_in <= "101010"; z_correct<="1110010010";
        when 174 => y_in <= "0110"; x_in <= "101010"; z_correct<="1101111100";
        when 175 => y_in <= "0111"; x_in <= "101010"; z_correct<="1101100110";
        when 176 => y_in <= "1000"; x_in <= "101011"; z_correct<="0010101000";
        when 177 => y_in <= "1001"; x_in <= "101011"; z_correct<="0010010011";
        when 178 => y_in <= "1010"; x_in <= "101011"; z_correct<="0001111110";
        when 179 => y_in <= "1011"; x_in <= "101011"; z_correct<="0001101001";
        when 180 => y_in <= "1100"; x_in <= "101011"; z_correct<="0001010100";
        when 181 => y_in <= "1101"; x_in <= "101011"; z_correct<="0000111111";
        when 182 => y_in <= "1110"; x_in <= "101011"; z_correct<="0000101010";
        when 183 => y_in <= "1111"; x_in <= "101011"; z_correct<="0000010101";
        when 184 => y_in <= "0000"; x_in <= "101011"; z_correct<="0000000000";
        when 185 => y_in <= "0001"; x_in <= "101011"; z_correct<="1111101011";
        when 186 => y_in <= "0010"; x_in <= "101011"; z_correct<="1111010110";
        when 187 => y_in <= "0011"; x_in <= "101011"; z_correct<="1111000001";
        when 188 => y_in <= "0100"; x_in <= "101011"; z_correct<="1110101100";
        when 189 => y_in <= "0101"; x_in <= "101011"; z_correct<="1110010111";
        when 190 => y_in <= "0110"; x_in <= "101011"; z_correct<="1110000010";
        when 191 => y_in <= "0111"; x_in <= "101011"; z_correct<="1101101101";
        when 192 => y_in <= "1000"; x_in <= "101100"; z_correct<="0010100000";
        when 193 => y_in <= "1001"; x_in <= "101100"; z_correct<="0010001100";
        when 194 => y_in <= "1010"; x_in <= "101100"; z_correct<="0001111000";
        when 195 => y_in <= "1011"; x_in <= "101100"; z_correct<="0001100100";
        when 196 => y_in <= "1100"; x_in <= "101100"; z_correct<="0001010000";
        when 197 => y_in <= "1101"; x_in <= "101100"; z_correct<="0000111100";
        when 198 => y_in <= "1110"; x_in <= "101100"; z_correct<="0000101000";
        when 199 => y_in <= "1111"; x_in <= "101100"; z_correct<="0000010100";
        when 200 => y_in <= "0000"; x_in <= "101100"; z_correct<="0000000000";
        when 201 => y_in <= "0001"; x_in <= "101100"; z_correct<="1111101100";
        when 202 => y_in <= "0010"; x_in <= "101100"; z_correct<="1111011000";
        when 203 => y_in <= "0011"; x_in <= "101100"; z_correct<="1111000100";
        when 204 => y_in <= "0100"; x_in <= "101100"; z_correct<="1110110000";
        when 205 => y_in <= "0101"; x_in <= "101100"; z_correct<="1110011100";
        when 206 => y_in <= "0110"; x_in <= "101100"; z_correct<="1110001000";
        when 207 => y_in <= "0111"; x_in <= "101100"; z_correct<="1101110100";
        when 208 => y_in <= "1000"; x_in <= "101101"; z_correct<="0010011000";
        when 209 => y_in <= "1001"; x_in <= "101101"; z_correct<="0010000101";
        when 210 => y_in <= "1010"; x_in <= "101101"; z_correct<="0001110010";
        when 211 => y_in <= "1011"; x_in <= "101101"; z_correct<="0001011111";
        when 212 => y_in <= "1100"; x_in <= "101101"; z_correct<="0001001100";
        when 213 => y_in <= "1101"; x_in <= "101101"; z_correct<="0000111001";
        when 214 => y_in <= "1110"; x_in <= "101101"; z_correct<="0000100110";
        when 215 => y_in <= "1111"; x_in <= "101101"; z_correct<="0000010011";
        when 216 => y_in <= "0000"; x_in <= "101101"; z_correct<="0000000000";
        when 217 => y_in <= "0001"; x_in <= "101101"; z_correct<="1111101101";
        when 218 => y_in <= "0010"; x_in <= "101101"; z_correct<="1111011010";
        when 219 => y_in <= "0011"; x_in <= "101101"; z_correct<="1111000111";
        when 220 => y_in <= "0100"; x_in <= "101101"; z_correct<="1110110100";
        when 221 => y_in <= "0101"; x_in <= "101101"; z_correct<="1110100001";
        when 222 => y_in <= "0110"; x_in <= "101101"; z_correct<="1110001110";
        when 223 => y_in <= "0111"; x_in <= "101101"; z_correct<="1101111011";
        when 224 => y_in <= "1000"; x_in <= "101110"; z_correct<="0010010000";
        when 225 => y_in <= "1001"; x_in <= "101110"; z_correct<="0001111110";
        when 226 => y_in <= "1010"; x_in <= "101110"; z_correct<="0001101100";
        when 227 => y_in <= "1011"; x_in <= "101110"; z_correct<="0001011010";
        when 228 => y_in <= "1100"; x_in <= "101110"; z_correct<="0001001000";
        when 229 => y_in <= "1101"; x_in <= "101110"; z_correct<="0000110110";
        when 230 => y_in <= "1110"; x_in <= "101110"; z_correct<="0000100100";
        when 231 => y_in <= "1111"; x_in <= "101110"; z_correct<="0000010010";
        when 232 => y_in <= "0000"; x_in <= "101110"; z_correct<="0000000000";
        when 233 => y_in <= "0001"; x_in <= "101110"; z_correct<="1111101110";
        when 234 => y_in <= "0010"; x_in <= "101110"; z_correct<="1111011100";
        when 235 => y_in <= "0011"; x_in <= "101110"; z_correct<="1111001010";
        when 236 => y_in <= "0100"; x_in <= "101110"; z_correct<="1110111000";
        when 237 => y_in <= "0101"; x_in <= "101110"; z_correct<="1110100110";
        when 238 => y_in <= "0110"; x_in <= "101110"; z_correct<="1110010100";
        when 239 => y_in <= "0111"; x_in <= "101110"; z_correct<="1110000010";
        when 240 => y_in <= "1000"; x_in <= "101111"; z_correct<="0010001000";
        when 241 => y_in <= "1001"; x_in <= "101111"; z_correct<="0001110111";
        when 242 => y_in <= "1010"; x_in <= "101111"; z_correct<="0001100110";
        when 243 => y_in <= "1011"; x_in <= "101111"; z_correct<="0001010101";
        when 244 => y_in <= "1100"; x_in <= "101111"; z_correct<="0001000100";
        when 245 => y_in <= "1101"; x_in <= "101111"; z_correct<="0000110011";
        when 246 => y_in <= "1110"; x_in <= "101111"; z_correct<="0000100010";
        when 247 => y_in <= "1111"; x_in <= "101111"; z_correct<="0000010001";
        when 248 => y_in <= "0000"; x_in <= "101111"; z_correct<="0000000000";
        when 249 => y_in <= "0001"; x_in <= "101111"; z_correct<="1111101111";
        when 250 => y_in <= "0010"; x_in <= "101111"; z_correct<="1111011110";
        when 251 => y_in <= "0011"; x_in <= "101111"; z_correct<="1111001101";
        when 252 => y_in <= "0100"; x_in <= "101111"; z_correct<="1110111100";
        when 253 => y_in <= "0101"; x_in <= "101111"; z_correct<="1110101011";
        when 254 => y_in <= "0110"; x_in <= "101111"; z_correct<="1110011010";
        when 255 => y_in <= "0111"; x_in <= "101111"; z_correct<="1110001001";
        when 256 => y_in <= "1000"; x_in <= "110000"; z_correct<="0010000000";
        when 257 => y_in <= "1001"; x_in <= "110000"; z_correct<="0001110000";
        when 258 => y_in <= "1010"; x_in <= "110000"; z_correct<="0001100000";
        when 259 => y_in <= "1011"; x_in <= "110000"; z_correct<="0001010000";
        when 260 => y_in <= "1100"; x_in <= "110000"; z_correct<="0001000000";
        when 261 => y_in <= "1101"; x_in <= "110000"; z_correct<="0000110000";
        when 262 => y_in <= "1110"; x_in <= "110000"; z_correct<="0000100000";
        when 263 => y_in <= "1111"; x_in <= "110000"; z_correct<="0000010000";
        when 264 => y_in <= "0000"; x_in <= "110000"; z_correct<="0000000000";
        when 265 => y_in <= "0001"; x_in <= "110000"; z_correct<="1111110000";
        when 266 => y_in <= "0010"; x_in <= "110000"; z_correct<="1111100000";
        when 267 => y_in <= "0011"; x_in <= "110000"; z_correct<="1111010000";
        when 268 => y_in <= "0100"; x_in <= "110000"; z_correct<="1111000000";
        when 269 => y_in <= "0101"; x_in <= "110000"; z_correct<="1110110000";
        when 270 => y_in <= "0110"; x_in <= "110000"; z_correct<="1110100000";
        when 271 => y_in <= "0111"; x_in <= "110000"; z_correct<="1110010000";
        when 272 => y_in <= "1000"; x_in <= "110001"; z_correct<="0001111000";
        when 273 => y_in <= "1001"; x_in <= "110001"; z_correct<="0001101001";
        when 274 => y_in <= "1010"; x_in <= "110001"; z_correct<="0001011010";
        when 275 => y_in <= "1011"; x_in <= "110001"; z_correct<="0001001011";
        when 276 => y_in <= "1100"; x_in <= "110001"; z_correct<="0000111100";
        when 277 => y_in <= "1101"; x_in <= "110001"; z_correct<="0000101101";
        when 278 => y_in <= "1110"; x_in <= "110001"; z_correct<="0000011110";
        when 279 => y_in <= "1111"; x_in <= "110001"; z_correct<="0000001111";
        when 280 => y_in <= "0000"; x_in <= "110001"; z_correct<="0000000000";
        when 281 => y_in <= "0001"; x_in <= "110001"; z_correct<="1111110001";
        when 282 => y_in <= "0010"; x_in <= "110001"; z_correct<="1111100010";
        when 283 => y_in <= "0011"; x_in <= "110001"; z_correct<="1111010011";
        when 284 => y_in <= "0100"; x_in <= "110001"; z_correct<="1111000100";
        when 285 => y_in <= "0101"; x_in <= "110001"; z_correct<="1110110101";
        when 286 => y_in <= "0110"; x_in <= "110001"; z_correct<="1110100110";
        when 287 => y_in <= "0111"; x_in <= "110001"; z_correct<="1110010111";
        when 288 => y_in <= "1000"; x_in <= "110010"; z_correct<="0001110000";
        when 289 => y_in <= "1001"; x_in <= "110010"; z_correct<="0001100010";
        when 290 => y_in <= "1010"; x_in <= "110010"; z_correct<="0001010100";
        when 291 => y_in <= "1011"; x_in <= "110010"; z_correct<="0001000110";
        when 292 => y_in <= "1100"; x_in <= "110010"; z_correct<="0000111000";
        when 293 => y_in <= "1101"; x_in <= "110010"; z_correct<="0000101010";
        when 294 => y_in <= "1110"; x_in <= "110010"; z_correct<="0000011100";
        when 295 => y_in <= "1111"; x_in <= "110010"; z_correct<="0000001110";
        when 296 => y_in <= "0000"; x_in <= "110010"; z_correct<="0000000000";
        when 297 => y_in <= "0001"; x_in <= "110010"; z_correct<="1111110010";
        when 298 => y_in <= "0010"; x_in <= "110010"; z_correct<="1111100100";
        when 299 => y_in <= "0011"; x_in <= "110010"; z_correct<="1111010110";
        when 300 => y_in <= "0100"; x_in <= "110010"; z_correct<="1111001000";
        when 301 => y_in <= "0101"; x_in <= "110010"; z_correct<="1110111010";
        when 302 => y_in <= "0110"; x_in <= "110010"; z_correct<="1110101100";
        when 303 => y_in <= "0111"; x_in <= "110010"; z_correct<="1110011110";
        when 304 => y_in <= "1000"; x_in <= "110011"; z_correct<="0001101000";
        when 305 => y_in <= "1001"; x_in <= "110011"; z_correct<="0001011011";
        when 306 => y_in <= "1010"; x_in <= "110011"; z_correct<="0001001110";
        when 307 => y_in <= "1011"; x_in <= "110011"; z_correct<="0001000001";
        when 308 => y_in <= "1100"; x_in <= "110011"; z_correct<="0000110100";
        when 309 => y_in <= "1101"; x_in <= "110011"; z_correct<="0000100111";
        when 310 => y_in <= "1110"; x_in <= "110011"; z_correct<="0000011010";
        when 311 => y_in <= "1111"; x_in <= "110011"; z_correct<="0000001101";
        when 312 => y_in <= "0000"; x_in <= "110011"; z_correct<="0000000000";
        when 313 => y_in <= "0001"; x_in <= "110011"; z_correct<="1111110011";
        when 314 => y_in <= "0010"; x_in <= "110011"; z_correct<="1111100110";
        when 315 => y_in <= "0011"; x_in <= "110011"; z_correct<="1111011001";
        when 316 => y_in <= "0100"; x_in <= "110011"; z_correct<="1111001100";
        when 317 => y_in <= "0101"; x_in <= "110011"; z_correct<="1110111111";
        when 318 => y_in <= "0110"; x_in <= "110011"; z_correct<="1110110010";
        when 319 => y_in <= "0111"; x_in <= "110011"; z_correct<="1110100101";
        when 320 => y_in <= "1000"; x_in <= "110100"; z_correct<="0001100000";
        when 321 => y_in <= "1001"; x_in <= "110100"; z_correct<="0001010100";
        when 322 => y_in <= "1010"; x_in <= "110100"; z_correct<="0001001000";
        when 323 => y_in <= "1011"; x_in <= "110100"; z_correct<="0000111100";
        when 324 => y_in <= "1100"; x_in <= "110100"; z_correct<="0000110000";
        when 325 => y_in <= "1101"; x_in <= "110100"; z_correct<="0000100100";
        when 326 => y_in <= "1110"; x_in <= "110100"; z_correct<="0000011000";
        when 327 => y_in <= "1111"; x_in <= "110100"; z_correct<="0000001100";
        when 328 => y_in <= "0000"; x_in <= "110100"; z_correct<="0000000000";
        when 329 => y_in <= "0001"; x_in <= "110100"; z_correct<="1111110100";
        when 330 => y_in <= "0010"; x_in <= "110100"; z_correct<="1111101000";
        when 331 => y_in <= "0011"; x_in <= "110100"; z_correct<="1111011100";
        when 332 => y_in <= "0100"; x_in <= "110100"; z_correct<="1111010000";
        when 333 => y_in <= "0101"; x_in <= "110100"; z_correct<="1111000100";
        when 334 => y_in <= "0110"; x_in <= "110100"; z_correct<="1110111000";
        when 335 => y_in <= "0111"; x_in <= "110100"; z_correct<="1110101100";
        when 336 => y_in <= "1000"; x_in <= "110101"; z_correct<="0001011000";
        when 337 => y_in <= "1001"; x_in <= "110101"; z_correct<="0001001101";
        when 338 => y_in <= "1010"; x_in <= "110101"; z_correct<="0001000010";
        when 339 => y_in <= "1011"; x_in <= "110101"; z_correct<="0000110111";
        when 340 => y_in <= "1100"; x_in <= "110101"; z_correct<="0000101100";
        when 341 => y_in <= "1101"; x_in <= "110101"; z_correct<="0000100001";
        when 342 => y_in <= "1110"; x_in <= "110101"; z_correct<="0000010110";
        when 343 => y_in <= "1111"; x_in <= "110101"; z_correct<="0000001011";
        when 344 => y_in <= "0000"; x_in <= "110101"; z_correct<="0000000000";
        when 345 => y_in <= "0001"; x_in <= "110101"; z_correct<="1111110101";
        when 346 => y_in <= "0010"; x_in <= "110101"; z_correct<="1111101010";
        when 347 => y_in <= "0011"; x_in <= "110101"; z_correct<="1111011111";
        when 348 => y_in <= "0100"; x_in <= "110101"; z_correct<="1111010100";
        when 349 => y_in <= "0101"; x_in <= "110101"; z_correct<="1111001001";
        when 350 => y_in <= "0110"; x_in <= "110101"; z_correct<="1110111110";
        when 351 => y_in <= "0111"; x_in <= "110101"; z_correct<="1110110011";
        when 352 => y_in <= "1000"; x_in <= "110110"; z_correct<="0001010000";
        when 353 => y_in <= "1001"; x_in <= "110110"; z_correct<="0001000110";
        when 354 => y_in <= "1010"; x_in <= "110110"; z_correct<="0000111100";
        when 355 => y_in <= "1011"; x_in <= "110110"; z_correct<="0000110010";
        when 356 => y_in <= "1100"; x_in <= "110110"; z_correct<="0000101000";
        when 357 => y_in <= "1101"; x_in <= "110110"; z_correct<="0000011110";
        when 358 => y_in <= "1110"; x_in <= "110110"; z_correct<="0000010100";
        when 359 => y_in <= "1111"; x_in <= "110110"; z_correct<="0000001010";
        when 360 => y_in <= "0000"; x_in <= "110110"; z_correct<="0000000000";
        when 361 => y_in <= "0001"; x_in <= "110110"; z_correct<="1111110110";
        when 362 => y_in <= "0010"; x_in <= "110110"; z_correct<="1111101100";
        when 363 => y_in <= "0011"; x_in <= "110110"; z_correct<="1111100010";
        when 364 => y_in <= "0100"; x_in <= "110110"; z_correct<="1111011000";
        when 365 => y_in <= "0101"; x_in <= "110110"; z_correct<="1111001110";
        when 366 => y_in <= "0110"; x_in <= "110110"; z_correct<="1111000100";
        when 367 => y_in <= "0111"; x_in <= "110110"; z_correct<="1110111010";
        when 368 => y_in <= "1000"; x_in <= "110111"; z_correct<="0001001000";
        when 369 => y_in <= "1001"; x_in <= "110111"; z_correct<="0000111111";
        when 370 => y_in <= "1010"; x_in <= "110111"; z_correct<="0000110110";
        when 371 => y_in <= "1011"; x_in <= "110111"; z_correct<="0000101101";
        when 372 => y_in <= "1100"; x_in <= "110111"; z_correct<="0000100100";
        when 373 => y_in <= "1101"; x_in <= "110111"; z_correct<="0000011011";
        when 374 => y_in <= "1110"; x_in <= "110111"; z_correct<="0000010010";
        when 375 => y_in <= "1111"; x_in <= "110111"; z_correct<="0000001001";
        when 376 => y_in <= "0000"; x_in <= "110111"; z_correct<="0000000000";
        when 377 => y_in <= "0001"; x_in <= "110111"; z_correct<="1111110111";
        when 378 => y_in <= "0010"; x_in <= "110111"; z_correct<="1111101110";
        when 379 => y_in <= "0011"; x_in <= "110111"; z_correct<="1111100101";
        when 380 => y_in <= "0100"; x_in <= "110111"; z_correct<="1111011100";
        when 381 => y_in <= "0101"; x_in <= "110111"; z_correct<="1111010011";
        when 382 => y_in <= "0110"; x_in <= "110111"; z_correct<="1111001010";
        when 383 => y_in <= "0111"; x_in <= "110111"; z_correct<="1111000001";
        when 384 => y_in <= "1000"; x_in <= "111000"; z_correct<="0001000000";
        when 385 => y_in <= "1001"; x_in <= "111000"; z_correct<="0000111000";
        when 386 => y_in <= "1010"; x_in <= "111000"; z_correct<="0000110000";
        when 387 => y_in <= "1011"; x_in <= "111000"; z_correct<="0000101000";
        when 388 => y_in <= "1100"; x_in <= "111000"; z_correct<="0000100000";
        when 389 => y_in <= "1101"; x_in <= "111000"; z_correct<="0000011000";
        when 390 => y_in <= "1110"; x_in <= "111000"; z_correct<="0000010000";
        when 391 => y_in <= "1111"; x_in <= "111000"; z_correct<="0000001000";
        when 392 => y_in <= "0000"; x_in <= "111000"; z_correct<="0000000000";
        when 393 => y_in <= "0001"; x_in <= "111000"; z_correct<="1111111000";
        when 394 => y_in <= "0010"; x_in <= "111000"; z_correct<="1111110000";
        when 395 => y_in <= "0011"; x_in <= "111000"; z_correct<="1111101000";
        when 396 => y_in <= "0100"; x_in <= "111000"; z_correct<="1111100000";
        when 397 => y_in <= "0101"; x_in <= "111000"; z_correct<="1111011000";
        when 398 => y_in <= "0110"; x_in <= "111000"; z_correct<="1111010000";
        when 399 => y_in <= "0111"; x_in <= "111000"; z_correct<="1111001000";
        when 400 => y_in <= "1000"; x_in <= "111001"; z_correct<="0000111000";
        when 401 => y_in <= "1001"; x_in <= "111001"; z_correct<="0000110001";
        when 402 => y_in <= "1010"; x_in <= "111001"; z_correct<="0000101010";
        when 403 => y_in <= "1011"; x_in <= "111001"; z_correct<="0000100011";
        when 404 => y_in <= "1100"; x_in <= "111001"; z_correct<="0000011100";
        when 405 => y_in <= "1101"; x_in <= "111001"; z_correct<="0000010101";
        when 406 => y_in <= "1110"; x_in <= "111001"; z_correct<="0000001110";
        when 407 => y_in <= "1111"; x_in <= "111001"; z_correct<="0000000111";
        when 408 => y_in <= "0000"; x_in <= "111001"; z_correct<="0000000000";
        when 409 => y_in <= "0001"; x_in <= "111001"; z_correct<="1111111001";
        when 410 => y_in <= "0010"; x_in <= "111001"; z_correct<="1111110010";
        when 411 => y_in <= "0011"; x_in <= "111001"; z_correct<="1111101011";
        when 412 => y_in <= "0100"; x_in <= "111001"; z_correct<="1111100100";
        when 413 => y_in <= "0101"; x_in <= "111001"; z_correct<="1111011101";
        when 414 => y_in <= "0110"; x_in <= "111001"; z_correct<="1111010110";
        when 415 => y_in <= "0111"; x_in <= "111001"; z_correct<="1111001111";
        when 416 => y_in <= "1000"; x_in <= "111010"; z_correct<="0000110000";
        when 417 => y_in <= "1001"; x_in <= "111010"; z_correct<="0000101010";
        when 418 => y_in <= "1010"; x_in <= "111010"; z_correct<="0000100100";
        when 419 => y_in <= "1011"; x_in <= "111010"; z_correct<="0000011110";
        when 420 => y_in <= "1100"; x_in <= "111010"; z_correct<="0000011000";
        when 421 => y_in <= "1101"; x_in <= "111010"; z_correct<="0000010010";
        when 422 => y_in <= "1110"; x_in <= "111010"; z_correct<="0000001100";
        when 423 => y_in <= "1111"; x_in <= "111010"; z_correct<="0000000110";
        when 424 => y_in <= "0000"; x_in <= "111010"; z_correct<="0000000000";
        when 425 => y_in <= "0001"; x_in <= "111010"; z_correct<="1111111010";
        when 426 => y_in <= "0010"; x_in <= "111010"; z_correct<="1111110100";
        when 427 => y_in <= "0011"; x_in <= "111010"; z_correct<="1111101110";
        when 428 => y_in <= "0100"; x_in <= "111010"; z_correct<="1111101000";
        when 429 => y_in <= "0101"; x_in <= "111010"; z_correct<="1111100010";
        when 430 => y_in <= "0110"; x_in <= "111010"; z_correct<="1111011100";
        when 431 => y_in <= "0111"; x_in <= "111010"; z_correct<="1111010110";
        when 432 => y_in <= "1000"; x_in <= "111011"; z_correct<="0000101000";
        when 433 => y_in <= "1001"; x_in <= "111011"; z_correct<="0000100011";
        when 434 => y_in <= "1010"; x_in <= "111011"; z_correct<="0000011110";
        when 435 => y_in <= "1011"; x_in <= "111011"; z_correct<="0000011001";
        when 436 => y_in <= "1100"; x_in <= "111011"; z_correct<="0000010100";
        when 437 => y_in <= "1101"; x_in <= "111011"; z_correct<="0000001111";
        when 438 => y_in <= "1110"; x_in <= "111011"; z_correct<="0000001010";
        when 439 => y_in <= "1111"; x_in <= "111011"; z_correct<="0000000101";
        when 440 => y_in <= "0000"; x_in <= "111011"; z_correct<="0000000000";
        when 441 => y_in <= "0001"; x_in <= "111011"; z_correct<="1111111011";
        when 442 => y_in <= "0010"; x_in <= "111011"; z_correct<="1111110110";
        when 443 => y_in <= "0011"; x_in <= "111011"; z_correct<="1111110001";
        when 444 => y_in <= "0100"; x_in <= "111011"; z_correct<="1111101100";
        when 445 => y_in <= "0101"; x_in <= "111011"; z_correct<="1111100111";
        when 446 => y_in <= "0110"; x_in <= "111011"; z_correct<="1111100010";
        when 447 => y_in <= "0111"; x_in <= "111011"; z_correct<="1111011101";
        when 448 => y_in <= "1000"; x_in <= "111100"; z_correct<="0000100000";
        when 449 => y_in <= "1001"; x_in <= "111100"; z_correct<="0000011100";
        when 450 => y_in <= "1010"; x_in <= "111100"; z_correct<="0000011000";
        when 451 => y_in <= "1011"; x_in <= "111100"; z_correct<="0000010100";
        when 452 => y_in <= "1100"; x_in <= "111100"; z_correct<="0000010000";
        when 453 => y_in <= "1101"; x_in <= "111100"; z_correct<="0000001100";
        when 454 => y_in <= "1110"; x_in <= "111100"; z_correct<="0000001000";
        when 455 => y_in <= "1111"; x_in <= "111100"; z_correct<="0000000100";
        when 456 => y_in <= "0000"; x_in <= "111100"; z_correct<="0000000000";
        when 457 => y_in <= "0001"; x_in <= "111100"; z_correct<="1111111100";
        when 458 => y_in <= "0010"; x_in <= "111100"; z_correct<="1111111000";
        when 459 => y_in <= "0011"; x_in <= "111100"; z_correct<="1111110100";
        when 460 => y_in <= "0100"; x_in <= "111100"; z_correct<="1111110000";
        when 461 => y_in <= "0101"; x_in <= "111100"; z_correct<="1111101100";
        when 462 => y_in <= "0110"; x_in <= "111100"; z_correct<="1111101000";
        when 463 => y_in <= "0111"; x_in <= "111100"; z_correct<="1111100100";
        when 464 => y_in <= "1000"; x_in <= "111101"; z_correct<="0000011000";
        when 465 => y_in <= "1001"; x_in <= "111101"; z_correct<="0000010101";
        when 466 => y_in <= "1010"; x_in <= "111101"; z_correct<="0000010010";
        when 467 => y_in <= "1011"; x_in <= "111101"; z_correct<="0000001111";
        when 468 => y_in <= "1100"; x_in <= "111101"; z_correct<="0000001100";
        when 469 => y_in <= "1101"; x_in <= "111101"; z_correct<="0000001001";
        when 470 => y_in <= "1110"; x_in <= "111101"; z_correct<="0000000110";
        when 471 => y_in <= "1111"; x_in <= "111101"; z_correct<="0000000011";
        when 472 => y_in <= "0000"; x_in <= "111101"; z_correct<="0000000000";
        when 473 => y_in <= "0001"; x_in <= "111101"; z_correct<="1111111101";
        when 474 => y_in <= "0010"; x_in <= "111101"; z_correct<="1111111010";
        when 475 => y_in <= "0011"; x_in <= "111101"; z_correct<="1111110111";
        when 476 => y_in <= "0100"; x_in <= "111101"; z_correct<="1111110100";
        when 477 => y_in <= "0101"; x_in <= "111101"; z_correct<="1111110001";
        when 478 => y_in <= "0110"; x_in <= "111101"; z_correct<="1111101110";
        when 479 => y_in <= "0111"; x_in <= "111101"; z_correct<="1111101011";
        when 480 => y_in <= "1000"; x_in <= "111110"; z_correct<="0000010000";
        when 481 => y_in <= "1001"; x_in <= "111110"; z_correct<="0000001110";
        when 482 => y_in <= "1010"; x_in <= "111110"; z_correct<="0000001100";
        when 483 => y_in <= "1011"; x_in <= "111110"; z_correct<="0000001010";
        when 484 => y_in <= "1100"; x_in <= "111110"; z_correct<="0000001000";
        when 485 => y_in <= "1101"; x_in <= "111110"; z_correct<="0000000110";
        when 486 => y_in <= "1110"; x_in <= "111110"; z_correct<="0000000100";
        when 487 => y_in <= "1111"; x_in <= "111110"; z_correct<="0000000010";
        when 488 => y_in <= "0000"; x_in <= "111110"; z_correct<="0000000000";
        when 489 => y_in <= "0001"; x_in <= "111110"; z_correct<="1111111110";
        when 490 => y_in <= "0010"; x_in <= "111110"; z_correct<="1111111100";
        when 491 => y_in <= "0011"; x_in <= "111110"; z_correct<="1111111010";
        when 492 => y_in <= "0100"; x_in <= "111110"; z_correct<="1111111000";
        when 493 => y_in <= "0101"; x_in <= "111110"; z_correct<="1111110110";
        when 494 => y_in <= "0110"; x_in <= "111110"; z_correct<="1111110100";
        when 495 => y_in <= "0111"; x_in <= "111110"; z_correct<="1111110010";
        when 496 => y_in <= "1000"; x_in <= "111111"; z_correct<="0000001000";
        when 497 => y_in <= "1001"; x_in <= "111111"; z_correct<="0000000111";
        when 498 => y_in <= "1010"; x_in <= "111111"; z_correct<="0000000110";
        when 499 => y_in <= "1011"; x_in <= "111111"; z_correct<="0000000101";
        when 500 => y_in <= "1100"; x_in <= "111111"; z_correct<="0000000100";
        when 501 => y_in <= "1101"; x_in <= "111111"; z_correct<="0000000011";
        when 502 => y_in <= "1110"; x_in <= "111111"; z_correct<="0000000010";
        when 503 => y_in <= "1111"; x_in <= "111111"; z_correct<="0000000001";
        when 504 => y_in <= "0000"; x_in <= "111111"; z_correct<="0000000000";
        when 505 => y_in <= "0001"; x_in <= "111111"; z_correct<="1111111111";
        when 506 => y_in <= "0010"; x_in <= "111111"; z_correct<="1111111110";
        when 507 => y_in <= "0011"; x_in <= "111111"; z_correct<="1111111101";
        when 508 => y_in <= "0100"; x_in <= "111111"; z_correct<="1111111100";
        when 509 => y_in <= "0101"; x_in <= "111111"; z_correct<="1111111011";
        when 510 => y_in <= "0110"; x_in <= "111111"; z_correct<="1111111010";
        when 511 => y_in <= "0111"; x_in <= "111111"; z_correct<="1111111001";
        when 512 => y_in <= "1000"; x_in <= "000000"; z_correct<="0000000000";
        when 513 => y_in <= "1001"; x_in <= "000000"; z_correct<="0000000000";
        when 514 => y_in <= "1010"; x_in <= "000000"; z_correct<="0000000000";
        when 515 => y_in <= "1011"; x_in <= "000000"; z_correct<="0000000000";
        when 516 => y_in <= "1100"; x_in <= "000000"; z_correct<="0000000000";
        when 517 => y_in <= "1101"; x_in <= "000000"; z_correct<="0000000000";
        when 518 => y_in <= "1110"; x_in <= "000000"; z_correct<="0000000000";
        when 519 => y_in <= "1111"; x_in <= "000000"; z_correct<="0000000000";
        when 520 => y_in <= "0000"; x_in <= "000000"; z_correct<="0000000000";
        when 521 => y_in <= "0001"; x_in <= "000000"; z_correct<="0000000000";
        when 522 => y_in <= "0010"; x_in <= "000000"; z_correct<="0000000000";
        when 523 => y_in <= "0011"; x_in <= "000000"; z_correct<="0000000000";
        when 524 => y_in <= "0100"; x_in <= "000000"; z_correct<="0000000000";
        when 525 => y_in <= "0101"; x_in <= "000000"; z_correct<="0000000000";
        when 526 => y_in <= "0110"; x_in <= "000000"; z_correct<="0000000000";
        when 527 => y_in <= "0111"; x_in <= "000000"; z_correct<="0000000000";
        when 528 => y_in <= "1000"; x_in <= "000001"; z_correct<="1111111000";
        when 529 => y_in <= "1001"; x_in <= "000001"; z_correct<="1111111001";
        when 530 => y_in <= "1010"; x_in <= "000001"; z_correct<="1111111010";
        when 531 => y_in <= "1011"; x_in <= "000001"; z_correct<="1111111011";
        when 532 => y_in <= "1100"; x_in <= "000001"; z_correct<="1111111100";
        when 533 => y_in <= "1101"; x_in <= "000001"; z_correct<="1111111101";
        when 534 => y_in <= "1110"; x_in <= "000001"; z_correct<="1111111110";
        when 535 => y_in <= "1111"; x_in <= "000001"; z_correct<="1111111111";
        when 536 => y_in <= "0000"; x_in <= "000001"; z_correct<="0000000000";
        when 537 => y_in <= "0001"; x_in <= "000001"; z_correct<="0000000001";
        when 538 => y_in <= "0010"; x_in <= "000001"; z_correct<="0000000010";
        when 539 => y_in <= "0011"; x_in <= "000001"; z_correct<="0000000011";
        when 540 => y_in <= "0100"; x_in <= "000001"; z_correct<="0000000100";
        when 541 => y_in <= "0101"; x_in <= "000001"; z_correct<="0000000101";
        when 542 => y_in <= "0110"; x_in <= "000001"; z_correct<="0000000110";
        when 543 => y_in <= "0111"; x_in <= "000001"; z_correct<="0000000111";
        when 544 => y_in <= "1000"; x_in <= "000010"; z_correct<="1111110000";
        when 545 => y_in <= "1001"; x_in <= "000010"; z_correct<="1111110010";
        when 546 => y_in <= "1010"; x_in <= "000010"; z_correct<="1111110100";
        when 547 => y_in <= "1011"; x_in <= "000010"; z_correct<="1111110110";
        when 548 => y_in <= "1100"; x_in <= "000010"; z_correct<="1111111000";
        when 549 => y_in <= "1101"; x_in <= "000010"; z_correct<="1111111010";
        when 550 => y_in <= "1110"; x_in <= "000010"; z_correct<="1111111100";
        when 551 => y_in <= "1111"; x_in <= "000010"; z_correct<="1111111110";
        when 552 => y_in <= "0000"; x_in <= "000010"; z_correct<="0000000000";
        when 553 => y_in <= "0001"; x_in <= "000010"; z_correct<="0000000010";
        when 554 => y_in <= "0010"; x_in <= "000010"; z_correct<="0000000100";
        when 555 => y_in <= "0011"; x_in <= "000010"; z_correct<="0000000110";
        when 556 => y_in <= "0100"; x_in <= "000010"; z_correct<="0000001000";
        when 557 => y_in <= "0101"; x_in <= "000010"; z_correct<="0000001010";
        when 558 => y_in <= "0110"; x_in <= "000010"; z_correct<="0000001100";
        when 559 => y_in <= "0111"; x_in <= "000010"; z_correct<="0000001110";
        when 560 => y_in <= "1000"; x_in <= "000011"; z_correct<="1111101000";
        when 561 => y_in <= "1001"; x_in <= "000011"; z_correct<="1111101011";
        when 562 => y_in <= "1010"; x_in <= "000011"; z_correct<="1111101110";
        when 563 => y_in <= "1011"; x_in <= "000011"; z_correct<="1111110001";
        when 564 => y_in <= "1100"; x_in <= "000011"; z_correct<="1111110100";
        when 565 => y_in <= "1101"; x_in <= "000011"; z_correct<="1111110111";
        when 566 => y_in <= "1110"; x_in <= "000011"; z_correct<="1111111010";
        when 567 => y_in <= "1111"; x_in <= "000011"; z_correct<="1111111101";
        when 568 => y_in <= "0000"; x_in <= "000011"; z_correct<="0000000000";
        when 569 => y_in <= "0001"; x_in <= "000011"; z_correct<="0000000011";
        when 570 => y_in <= "0010"; x_in <= "000011"; z_correct<="0000000110";
        when 571 => y_in <= "0011"; x_in <= "000011"; z_correct<="0000001001";
        when 572 => y_in <= "0100"; x_in <= "000011"; z_correct<="0000001100";
        when 573 => y_in <= "0101"; x_in <= "000011"; z_correct<="0000001111";
        when 574 => y_in <= "0110"; x_in <= "000011"; z_correct<="0000010010";
        when 575 => y_in <= "0111"; x_in <= "000011"; z_correct<="0000010101";
        when 576 => y_in <= "1000"; x_in <= "000100"; z_correct<="1111100000";
        when 577 => y_in <= "1001"; x_in <= "000100"; z_correct<="1111100100";
        when 578 => y_in <= "1010"; x_in <= "000100"; z_correct<="1111101000";
        when 579 => y_in <= "1011"; x_in <= "000100"; z_correct<="1111101100";
        when 580 => y_in <= "1100"; x_in <= "000100"; z_correct<="1111110000";
        when 581 => y_in <= "1101"; x_in <= "000100"; z_correct<="1111110100";
        when 582 => y_in <= "1110"; x_in <= "000100"; z_correct<="1111111000";
        when 583 => y_in <= "1111"; x_in <= "000100"; z_correct<="1111111100";
        when 584 => y_in <= "0000"; x_in <= "000100"; z_correct<="0000000000";
        when 585 => y_in <= "0001"; x_in <= "000100"; z_correct<="0000000100";
        when 586 => y_in <= "0010"; x_in <= "000100"; z_correct<="0000001000";
        when 587 => y_in <= "0011"; x_in <= "000100"; z_correct<="0000001100";
        when 588 => y_in <= "0100"; x_in <= "000100"; z_correct<="0000010000";
        when 589 => y_in <= "0101"; x_in <= "000100"; z_correct<="0000010100";
        when 590 => y_in <= "0110"; x_in <= "000100"; z_correct<="0000011000";
        when 591 => y_in <= "0111"; x_in <= "000100"; z_correct<="0000011100";
        when 592 => y_in <= "1000"; x_in <= "000101"; z_correct<="1111011000";
        when 593 => y_in <= "1001"; x_in <= "000101"; z_correct<="1111011101";
        when 594 => y_in <= "1010"; x_in <= "000101"; z_correct<="1111100010";
        when 595 => y_in <= "1011"; x_in <= "000101"; z_correct<="1111100111";
        when 596 => y_in <= "1100"; x_in <= "000101"; z_correct<="1111101100";
        when 597 => y_in <= "1101"; x_in <= "000101"; z_correct<="1111110001";
        when 598 => y_in <= "1110"; x_in <= "000101"; z_correct<="1111110110";
        when 599 => y_in <= "1111"; x_in <= "000101"; z_correct<="1111111011";
        when 600 => y_in <= "0000"; x_in <= "000101"; z_correct<="0000000000";
        when 601 => y_in <= "0001"; x_in <= "000101"; z_correct<="0000000101";
        when 602 => y_in <= "0010"; x_in <= "000101"; z_correct<="0000001010";
        when 603 => y_in <= "0011"; x_in <= "000101"; z_correct<="0000001111";
        when 604 => y_in <= "0100"; x_in <= "000101"; z_correct<="0000010100";
        when 605 => y_in <= "0101"; x_in <= "000101"; z_correct<="0000011001";
        when 606 => y_in <= "0110"; x_in <= "000101"; z_correct<="0000011110";
        when 607 => y_in <= "0111"; x_in <= "000101"; z_correct<="0000100011";
        when 608 => y_in <= "1000"; x_in <= "000110"; z_correct<="1111010000";
        when 609 => y_in <= "1001"; x_in <= "000110"; z_correct<="1111010110";
        when 610 => y_in <= "1010"; x_in <= "000110"; z_correct<="1111011100";
        when 611 => y_in <= "1011"; x_in <= "000110"; z_correct<="1111100010";
        when 612 => y_in <= "1100"; x_in <= "000110"; z_correct<="1111101000";
        when 613 => y_in <= "1101"; x_in <= "000110"; z_correct<="1111101110";
        when 614 => y_in <= "1110"; x_in <= "000110"; z_correct<="1111110100";
        when 615 => y_in <= "1111"; x_in <= "000110"; z_correct<="1111111010";
        when 616 => y_in <= "0000"; x_in <= "000110"; z_correct<="0000000000";
        when 617 => y_in <= "0001"; x_in <= "000110"; z_correct<="0000000110";
        when 618 => y_in <= "0010"; x_in <= "000110"; z_correct<="0000001100";
        when 619 => y_in <= "0011"; x_in <= "000110"; z_correct<="0000010010";
        when 620 => y_in <= "0100"; x_in <= "000110"; z_correct<="0000011000";
        when 621 => y_in <= "0101"; x_in <= "000110"; z_correct<="0000011110";
        when 622 => y_in <= "0110"; x_in <= "000110"; z_correct<="0000100100";
        when 623 => y_in <= "0111"; x_in <= "000110"; z_correct<="0000101010";
        when 624 => y_in <= "1000"; x_in <= "000111"; z_correct<="1111001000";
        when 625 => y_in <= "1001"; x_in <= "000111"; z_correct<="1111001111";
        when 626 => y_in <= "1010"; x_in <= "000111"; z_correct<="1111010110";
        when 627 => y_in <= "1011"; x_in <= "000111"; z_correct<="1111011101";
        when 628 => y_in <= "1100"; x_in <= "000111"; z_correct<="1111100100";
        when 629 => y_in <= "1101"; x_in <= "000111"; z_correct<="1111101011";
        when 630 => y_in <= "1110"; x_in <= "000111"; z_correct<="1111110010";
        when 631 => y_in <= "1111"; x_in <= "000111"; z_correct<="1111111001";
        when 632 => y_in <= "0000"; x_in <= "000111"; z_correct<="0000000000";
        when 633 => y_in <= "0001"; x_in <= "000111"; z_correct<="0000000111";
        when 634 => y_in <= "0010"; x_in <= "000111"; z_correct<="0000001110";
        when 635 => y_in <= "0011"; x_in <= "000111"; z_correct<="0000010101";
        when 636 => y_in <= "0100"; x_in <= "000111"; z_correct<="0000011100";
        when 637 => y_in <= "0101"; x_in <= "000111"; z_correct<="0000100011";
        when 638 => y_in <= "0110"; x_in <= "000111"; z_correct<="0000101010";
        when 639 => y_in <= "0111"; x_in <= "000111"; z_correct<="0000110001";
        when 640 => y_in <= "1000"; x_in <= "001000"; z_correct<="1111000000";
        when 641 => y_in <= "1001"; x_in <= "001000"; z_correct<="1111001000";
        when 642 => y_in <= "1010"; x_in <= "001000"; z_correct<="1111010000";
        when 643 => y_in <= "1011"; x_in <= "001000"; z_correct<="1111011000";
        when 644 => y_in <= "1100"; x_in <= "001000"; z_correct<="1111100000";
        when 645 => y_in <= "1101"; x_in <= "001000"; z_correct<="1111101000";
        when 646 => y_in <= "1110"; x_in <= "001000"; z_correct<="1111110000";
        when 647 => y_in <= "1111"; x_in <= "001000"; z_correct<="1111111000";
        when 648 => y_in <= "0000"; x_in <= "001000"; z_correct<="0000000000";
        when 649 => y_in <= "0001"; x_in <= "001000"; z_correct<="0000001000";
        when 650 => y_in <= "0010"; x_in <= "001000"; z_correct<="0000010000";
        when 651 => y_in <= "0011"; x_in <= "001000"; z_correct<="0000011000";
        when 652 => y_in <= "0100"; x_in <= "001000"; z_correct<="0000100000";
        when 653 => y_in <= "0101"; x_in <= "001000"; z_correct<="0000101000";
        when 654 => y_in <= "0110"; x_in <= "001000"; z_correct<="0000110000";
        when 655 => y_in <= "0111"; x_in <= "001000"; z_correct<="0000111000";
        when 656 => y_in <= "1000"; x_in <= "001001"; z_correct<="1110111000";
        when 657 => y_in <= "1001"; x_in <= "001001"; z_correct<="1111000001";
        when 658 => y_in <= "1010"; x_in <= "001001"; z_correct<="1111001010";
        when 659 => y_in <= "1011"; x_in <= "001001"; z_correct<="1111010011";
        when 660 => y_in <= "1100"; x_in <= "001001"; z_correct<="1111011100";
        when 661 => y_in <= "1101"; x_in <= "001001"; z_correct<="1111100101";
        when 662 => y_in <= "1110"; x_in <= "001001"; z_correct<="1111101110";
        when 663 => y_in <= "1111"; x_in <= "001001"; z_correct<="1111110111";
        when 664 => y_in <= "0000"; x_in <= "001001"; z_correct<="0000000000";
        when 665 => y_in <= "0001"; x_in <= "001001"; z_correct<="0000001001";
        when 666 => y_in <= "0010"; x_in <= "001001"; z_correct<="0000010010";
        when 667 => y_in <= "0011"; x_in <= "001001"; z_correct<="0000011011";
        when 668 => y_in <= "0100"; x_in <= "001001"; z_correct<="0000100100";
        when 669 => y_in <= "0101"; x_in <= "001001"; z_correct<="0000101101";
        when 670 => y_in <= "0110"; x_in <= "001001"; z_correct<="0000110110";
        when 671 => y_in <= "0111"; x_in <= "001001"; z_correct<="0000111111";
        when 672 => y_in <= "1000"; x_in <= "001010"; z_correct<="1110110000";
        when 673 => y_in <= "1001"; x_in <= "001010"; z_correct<="1110111010";
        when 674 => y_in <= "1010"; x_in <= "001010"; z_correct<="1111000100";
        when 675 => y_in <= "1011"; x_in <= "001010"; z_correct<="1111001110";
        when 676 => y_in <= "1100"; x_in <= "001010"; z_correct<="1111011000";
        when 677 => y_in <= "1101"; x_in <= "001010"; z_correct<="1111100010";
        when 678 => y_in <= "1110"; x_in <= "001010"; z_correct<="1111101100";
        when 679 => y_in <= "1111"; x_in <= "001010"; z_correct<="1111110110";
        when 680 => y_in <= "0000"; x_in <= "001010"; z_correct<="0000000000";
        when 681 => y_in <= "0001"; x_in <= "001010"; z_correct<="0000001010";
        when 682 => y_in <= "0010"; x_in <= "001010"; z_correct<="0000010100";
        when 683 => y_in <= "0011"; x_in <= "001010"; z_correct<="0000011110";
        when 684 => y_in <= "0100"; x_in <= "001010"; z_correct<="0000101000";
        when 685 => y_in <= "0101"; x_in <= "001010"; z_correct<="0000110010";
        when 686 => y_in <= "0110"; x_in <= "001010"; z_correct<="0000111100";
        when 687 => y_in <= "0111"; x_in <= "001010"; z_correct<="0001000110";
        when 688 => y_in <= "1000"; x_in <= "001011"; z_correct<="1110101000";
        when 689 => y_in <= "1001"; x_in <= "001011"; z_correct<="1110110011";
        when 690 => y_in <= "1010"; x_in <= "001011"; z_correct<="1110111110";
        when 691 => y_in <= "1011"; x_in <= "001011"; z_correct<="1111001001";
        when 692 => y_in <= "1100"; x_in <= "001011"; z_correct<="1111010100";
        when 693 => y_in <= "1101"; x_in <= "001011"; z_correct<="1111011111";
        when 694 => y_in <= "1110"; x_in <= "001011"; z_correct<="1111101010";
        when 695 => y_in <= "1111"; x_in <= "001011"; z_correct<="1111110101";
        when 696 => y_in <= "0000"; x_in <= "001011"; z_correct<="0000000000";
        when 697 => y_in <= "0001"; x_in <= "001011"; z_correct<="0000001011";
        when 698 => y_in <= "0010"; x_in <= "001011"; z_correct<="0000010110";
        when 699 => y_in <= "0011"; x_in <= "001011"; z_correct<="0000100001";
        when 700 => y_in <= "0100"; x_in <= "001011"; z_correct<="0000101100";
        when 701 => y_in <= "0101"; x_in <= "001011"; z_correct<="0000110111";
        when 702 => y_in <= "0110"; x_in <= "001011"; z_correct<="0001000010";
        when 703 => y_in <= "0111"; x_in <= "001011"; z_correct<="0001001101";
        when 704 => y_in <= "1000"; x_in <= "001100"; z_correct<="1110100000";
        when 705 => y_in <= "1001"; x_in <= "001100"; z_correct<="1110101100";
        when 706 => y_in <= "1010"; x_in <= "001100"; z_correct<="1110111000";
        when 707 => y_in <= "1011"; x_in <= "001100"; z_correct<="1111000100";
        when 708 => y_in <= "1100"; x_in <= "001100"; z_correct<="1111010000";
        when 709 => y_in <= "1101"; x_in <= "001100"; z_correct<="1111011100";
        when 710 => y_in <= "1110"; x_in <= "001100"; z_correct<="1111101000";
        when 711 => y_in <= "1111"; x_in <= "001100"; z_correct<="1111110100";
        when 712 => y_in <= "0000"; x_in <= "001100"; z_correct<="0000000000";
        when 713 => y_in <= "0001"; x_in <= "001100"; z_correct<="0000001100";
        when 714 => y_in <= "0010"; x_in <= "001100"; z_correct<="0000011000";
        when 715 => y_in <= "0011"; x_in <= "001100"; z_correct<="0000100100";
        when 716 => y_in <= "0100"; x_in <= "001100"; z_correct<="0000110000";
        when 717 => y_in <= "0101"; x_in <= "001100"; z_correct<="0000111100";
        when 718 => y_in <= "0110"; x_in <= "001100"; z_correct<="0001001000";
        when 719 => y_in <= "0111"; x_in <= "001100"; z_correct<="0001010100";
        when 720 => y_in <= "1000"; x_in <= "001101"; z_correct<="1110011000";
        when 721 => y_in <= "1001"; x_in <= "001101"; z_correct<="1110100101";
        when 722 => y_in <= "1010"; x_in <= "001101"; z_correct<="1110110010";
        when 723 => y_in <= "1011"; x_in <= "001101"; z_correct<="1110111111";
        when 724 => y_in <= "1100"; x_in <= "001101"; z_correct<="1111001100";
        when 725 => y_in <= "1101"; x_in <= "001101"; z_correct<="1111011001";
        when 726 => y_in <= "1110"; x_in <= "001101"; z_correct<="1111100110";
        when 727 => y_in <= "1111"; x_in <= "001101"; z_correct<="1111110011";
        when 728 => y_in <= "0000"; x_in <= "001101"; z_correct<="0000000000";
        when 729 => y_in <= "0001"; x_in <= "001101"; z_correct<="0000001101";
        when 730 => y_in <= "0010"; x_in <= "001101"; z_correct<="0000011010";
        when 731 => y_in <= "0011"; x_in <= "001101"; z_correct<="0000100111";
        when 732 => y_in <= "0100"; x_in <= "001101"; z_correct<="0000110100";
        when 733 => y_in <= "0101"; x_in <= "001101"; z_correct<="0001000001";
        when 734 => y_in <= "0110"; x_in <= "001101"; z_correct<="0001001110";
        when 735 => y_in <= "0111"; x_in <= "001101"; z_correct<="0001011011";
        when 736 => y_in <= "1000"; x_in <= "001110"; z_correct<="1110010000";
        when 737 => y_in <= "1001"; x_in <= "001110"; z_correct<="1110011110";
        when 738 => y_in <= "1010"; x_in <= "001110"; z_correct<="1110101100";
        when 739 => y_in <= "1011"; x_in <= "001110"; z_correct<="1110111010";
        when 740 => y_in <= "1100"; x_in <= "001110"; z_correct<="1111001000";
        when 741 => y_in <= "1101"; x_in <= "001110"; z_correct<="1111010110";
        when 742 => y_in <= "1110"; x_in <= "001110"; z_correct<="1111100100";
        when 743 => y_in <= "1111"; x_in <= "001110"; z_correct<="1111110010";
        when 744 => y_in <= "0000"; x_in <= "001110"; z_correct<="0000000000";
        when 745 => y_in <= "0001"; x_in <= "001110"; z_correct<="0000001110";
        when 746 => y_in <= "0010"; x_in <= "001110"; z_correct<="0000011100";
        when 747 => y_in <= "0011"; x_in <= "001110"; z_correct<="0000101010";
        when 748 => y_in <= "0100"; x_in <= "001110"; z_correct<="0000111000";
        when 749 => y_in <= "0101"; x_in <= "001110"; z_correct<="0001000110";
        when 750 => y_in <= "0110"; x_in <= "001110"; z_correct<="0001010100";
        when 751 => y_in <= "0111"; x_in <= "001110"; z_correct<="0001100010";
        when 752 => y_in <= "1000"; x_in <= "001111"; z_correct<="1110001000";
        when 753 => y_in <= "1001"; x_in <= "001111"; z_correct<="1110010111";
        when 754 => y_in <= "1010"; x_in <= "001111"; z_correct<="1110100110";
        when 755 => y_in <= "1011"; x_in <= "001111"; z_correct<="1110110101";
        when 756 => y_in <= "1100"; x_in <= "001111"; z_correct<="1111000100";
        when 757 => y_in <= "1101"; x_in <= "001111"; z_correct<="1111010011";
        when 758 => y_in <= "1110"; x_in <= "001111"; z_correct<="1111100010";
        when 759 => y_in <= "1111"; x_in <= "001111"; z_correct<="1111110001";
        when 760 => y_in <= "0000"; x_in <= "001111"; z_correct<="0000000000";
        when 761 => y_in <= "0001"; x_in <= "001111"; z_correct<="0000001111";
        when 762 => y_in <= "0010"; x_in <= "001111"; z_correct<="0000011110";
        when 763 => y_in <= "0011"; x_in <= "001111"; z_correct<="0000101101";
        when 764 => y_in <= "0100"; x_in <= "001111"; z_correct<="0000111100";
        when 765 => y_in <= "0101"; x_in <= "001111"; z_correct<="0001001011";
        when 766 => y_in <= "0110"; x_in <= "001111"; z_correct<="0001011010";
        when 767 => y_in <= "0111"; x_in <= "001111"; z_correct<="0001101001";
        when 768 => y_in <= "1000"; x_in <= "010000"; z_correct<="1110000000";
        when 769 => y_in <= "1001"; x_in <= "010000"; z_correct<="1110010000";
        when 770 => y_in <= "1010"; x_in <= "010000"; z_correct<="1110100000";
        when 771 => y_in <= "1011"; x_in <= "010000"; z_correct<="1110110000";
        when 772 => y_in <= "1100"; x_in <= "010000"; z_correct<="1111000000";
        when 773 => y_in <= "1101"; x_in <= "010000"; z_correct<="1111010000";
        when 774 => y_in <= "1110"; x_in <= "010000"; z_correct<="1111100000";
        when 775 => y_in <= "1111"; x_in <= "010000"; z_correct<="1111110000";
        when 776 => y_in <= "0000"; x_in <= "010000"; z_correct<="0000000000";
        when 777 => y_in <= "0001"; x_in <= "010000"; z_correct<="0000010000";
        when 778 => y_in <= "0010"; x_in <= "010000"; z_correct<="0000100000";
        when 779 => y_in <= "0011"; x_in <= "010000"; z_correct<="0000110000";
        when 780 => y_in <= "0100"; x_in <= "010000"; z_correct<="0001000000";
        when 781 => y_in <= "0101"; x_in <= "010000"; z_correct<="0001010000";
        when 782 => y_in <= "0110"; x_in <= "010000"; z_correct<="0001100000";
        when 783 => y_in <= "0111"; x_in <= "010000"; z_correct<="0001110000";
        when 784 => y_in <= "1000"; x_in <= "010001"; z_correct<="1101111000";
        when 785 => y_in <= "1001"; x_in <= "010001"; z_correct<="1110001001";
        when 786 => y_in <= "1010"; x_in <= "010001"; z_correct<="1110011010";
        when 787 => y_in <= "1011"; x_in <= "010001"; z_correct<="1110101011";
        when 788 => y_in <= "1100"; x_in <= "010001"; z_correct<="1110111100";
        when 789 => y_in <= "1101"; x_in <= "010001"; z_correct<="1111001101";
        when 790 => y_in <= "1110"; x_in <= "010001"; z_correct<="1111011110";
        when 791 => y_in <= "1111"; x_in <= "010001"; z_correct<="1111101111";
        when 792 => y_in <= "0000"; x_in <= "010001"; z_correct<="0000000000";
        when 793 => y_in <= "0001"; x_in <= "010001"; z_correct<="0000010001";
        when 794 => y_in <= "0010"; x_in <= "010001"; z_correct<="0000100010";
        when 795 => y_in <= "0011"; x_in <= "010001"; z_correct<="0000110011";
        when 796 => y_in <= "0100"; x_in <= "010001"; z_correct<="0001000100";
        when 797 => y_in <= "0101"; x_in <= "010001"; z_correct<="0001010101";
        when 798 => y_in <= "0110"; x_in <= "010001"; z_correct<="0001100110";
        when 799 => y_in <= "0111"; x_in <= "010001"; z_correct<="0001110111";
        when 800 => y_in <= "1000"; x_in <= "010010"; z_correct<="1101110000";
        when 801 => y_in <= "1001"; x_in <= "010010"; z_correct<="1110000010";
        when 802 => y_in <= "1010"; x_in <= "010010"; z_correct<="1110010100";
        when 803 => y_in <= "1011"; x_in <= "010010"; z_correct<="1110100110";
        when 804 => y_in <= "1100"; x_in <= "010010"; z_correct<="1110111000";
        when 805 => y_in <= "1101"; x_in <= "010010"; z_correct<="1111001010";
        when 806 => y_in <= "1110"; x_in <= "010010"; z_correct<="1111011100";
        when 807 => y_in <= "1111"; x_in <= "010010"; z_correct<="1111101110";
        when 808 => y_in <= "0000"; x_in <= "010010"; z_correct<="0000000000";
        when 809 => y_in <= "0001"; x_in <= "010010"; z_correct<="0000010010";
        when 810 => y_in <= "0010"; x_in <= "010010"; z_correct<="0000100100";
        when 811 => y_in <= "0011"; x_in <= "010010"; z_correct<="0000110110";
        when 812 => y_in <= "0100"; x_in <= "010010"; z_correct<="0001001000";
        when 813 => y_in <= "0101"; x_in <= "010010"; z_correct<="0001011010";
        when 814 => y_in <= "0110"; x_in <= "010010"; z_correct<="0001101100";
        when 815 => y_in <= "0111"; x_in <= "010010"; z_correct<="0001111110";
        when 816 => y_in <= "1000"; x_in <= "010011"; z_correct<="1101101000";
        when 817 => y_in <= "1001"; x_in <= "010011"; z_correct<="1101111011";
        when 818 => y_in <= "1010"; x_in <= "010011"; z_correct<="1110001110";
        when 819 => y_in <= "1011"; x_in <= "010011"; z_correct<="1110100001";
        when 820 => y_in <= "1100"; x_in <= "010011"; z_correct<="1110110100";
        when 821 => y_in <= "1101"; x_in <= "010011"; z_correct<="1111000111";
        when 822 => y_in <= "1110"; x_in <= "010011"; z_correct<="1111011010";
        when 823 => y_in <= "1111"; x_in <= "010011"; z_correct<="1111101101";
        when 824 => y_in <= "0000"; x_in <= "010011"; z_correct<="0000000000";
        when 825 => y_in <= "0001"; x_in <= "010011"; z_correct<="0000010011";
        when 826 => y_in <= "0010"; x_in <= "010011"; z_correct<="0000100110";
        when 827 => y_in <= "0011"; x_in <= "010011"; z_correct<="0000111001";
        when 828 => y_in <= "0100"; x_in <= "010011"; z_correct<="0001001100";
        when 829 => y_in <= "0101"; x_in <= "010011"; z_correct<="0001011111";
        when 830 => y_in <= "0110"; x_in <= "010011"; z_correct<="0001110010";
        when 831 => y_in <= "0111"; x_in <= "010011"; z_correct<="0010000101";
        when 832 => y_in <= "1000"; x_in <= "010100"; z_correct<="1101100000";
        when 833 => y_in <= "1001"; x_in <= "010100"; z_correct<="1101110100";
        when 834 => y_in <= "1010"; x_in <= "010100"; z_correct<="1110001000";
        when 835 => y_in <= "1011"; x_in <= "010100"; z_correct<="1110011100";
        when 836 => y_in <= "1100"; x_in <= "010100"; z_correct<="1110110000";
        when 837 => y_in <= "1101"; x_in <= "010100"; z_correct<="1111000100";
        when 838 => y_in <= "1110"; x_in <= "010100"; z_correct<="1111011000";
        when 839 => y_in <= "1111"; x_in <= "010100"; z_correct<="1111101100";
        when 840 => y_in <= "0000"; x_in <= "010100"; z_correct<="0000000000";
        when 841 => y_in <= "0001"; x_in <= "010100"; z_correct<="0000010100";
        when 842 => y_in <= "0010"; x_in <= "010100"; z_correct<="0000101000";
        when 843 => y_in <= "0011"; x_in <= "010100"; z_correct<="0000111100";
        when 844 => y_in <= "0100"; x_in <= "010100"; z_correct<="0001010000";
        when 845 => y_in <= "0101"; x_in <= "010100"; z_correct<="0001100100";
        when 846 => y_in <= "0110"; x_in <= "010100"; z_correct<="0001111000";
        when 847 => y_in <= "0111"; x_in <= "010100"; z_correct<="0010001100";
        when 848 => y_in <= "1000"; x_in <= "010101"; z_correct<="1101011000";
        when 849 => y_in <= "1001"; x_in <= "010101"; z_correct<="1101101101";
        when 850 => y_in <= "1010"; x_in <= "010101"; z_correct<="1110000010";
        when 851 => y_in <= "1011"; x_in <= "010101"; z_correct<="1110010111";
        when 852 => y_in <= "1100"; x_in <= "010101"; z_correct<="1110101100";
        when 853 => y_in <= "1101"; x_in <= "010101"; z_correct<="1111000001";
        when 854 => y_in <= "1110"; x_in <= "010101"; z_correct<="1111010110";
        when 855 => y_in <= "1111"; x_in <= "010101"; z_correct<="1111101011";
        when 856 => y_in <= "0000"; x_in <= "010101"; z_correct<="0000000000";
        when 857 => y_in <= "0001"; x_in <= "010101"; z_correct<="0000010101";
        when 858 => y_in <= "0010"; x_in <= "010101"; z_correct<="0000101010";
        when 859 => y_in <= "0011"; x_in <= "010101"; z_correct<="0000111111";
        when 860 => y_in <= "0100"; x_in <= "010101"; z_correct<="0001010100";
        when 861 => y_in <= "0101"; x_in <= "010101"; z_correct<="0001101001";
        when 862 => y_in <= "0110"; x_in <= "010101"; z_correct<="0001111110";
        when 863 => y_in <= "0111"; x_in <= "010101"; z_correct<="0010010011";
        when 864 => y_in <= "1000"; x_in <= "010110"; z_correct<="1101010000";
        when 865 => y_in <= "1001"; x_in <= "010110"; z_correct<="1101100110";
        when 866 => y_in <= "1010"; x_in <= "010110"; z_correct<="1101111100";
        when 867 => y_in <= "1011"; x_in <= "010110"; z_correct<="1110010010";
        when 868 => y_in <= "1100"; x_in <= "010110"; z_correct<="1110101000";
        when 869 => y_in <= "1101"; x_in <= "010110"; z_correct<="1110111110";
        when 870 => y_in <= "1110"; x_in <= "010110"; z_correct<="1111010100";
        when 871 => y_in <= "1111"; x_in <= "010110"; z_correct<="1111101010";
        when 872 => y_in <= "0000"; x_in <= "010110"; z_correct<="0000000000";
        when 873 => y_in <= "0001"; x_in <= "010110"; z_correct<="0000010110";
        when 874 => y_in <= "0010"; x_in <= "010110"; z_correct<="0000101100";
        when 875 => y_in <= "0011"; x_in <= "010110"; z_correct<="0001000010";
        when 876 => y_in <= "0100"; x_in <= "010110"; z_correct<="0001011000";
        when 877 => y_in <= "0101"; x_in <= "010110"; z_correct<="0001101110";
        when 878 => y_in <= "0110"; x_in <= "010110"; z_correct<="0010000100";
        when 879 => y_in <= "0111"; x_in <= "010110"; z_correct<="0010011010";
        when 880 => y_in <= "1000"; x_in <= "010111"; z_correct<="1101001000";
        when 881 => y_in <= "1001"; x_in <= "010111"; z_correct<="1101011111";
        when 882 => y_in <= "1010"; x_in <= "010111"; z_correct<="1101110110";
        when 883 => y_in <= "1011"; x_in <= "010111"; z_correct<="1110001101";
        when 884 => y_in <= "1100"; x_in <= "010111"; z_correct<="1110100100";
        when 885 => y_in <= "1101"; x_in <= "010111"; z_correct<="1110111011";
        when 886 => y_in <= "1110"; x_in <= "010111"; z_correct<="1111010010";
        when 887 => y_in <= "1111"; x_in <= "010111"; z_correct<="1111101001";
        when 888 => y_in <= "0000"; x_in <= "010111"; z_correct<="0000000000";
        when 889 => y_in <= "0001"; x_in <= "010111"; z_correct<="0000010111";
        when 890 => y_in <= "0010"; x_in <= "010111"; z_correct<="0000101110";
        when 891 => y_in <= "0011"; x_in <= "010111"; z_correct<="0001000101";
        when 892 => y_in <= "0100"; x_in <= "010111"; z_correct<="0001011100";
        when 893 => y_in <= "0101"; x_in <= "010111"; z_correct<="0001110011";
        when 894 => y_in <= "0110"; x_in <= "010111"; z_correct<="0010001010";
        when 895 => y_in <= "0111"; x_in <= "010111"; z_correct<="0010100001";
        when 896 => y_in <= "1000"; x_in <= "011000"; z_correct<="1101000000";
        when 897 => y_in <= "1001"; x_in <= "011000"; z_correct<="1101011000";
        when 898 => y_in <= "1010"; x_in <= "011000"; z_correct<="1101110000";
        when 899 => y_in <= "1011"; x_in <= "011000"; z_correct<="1110001000";
        when 900 => y_in <= "1100"; x_in <= "011000"; z_correct<="1110100000";
        when 901 => y_in <= "1101"; x_in <= "011000"; z_correct<="1110111000";
        when 902 => y_in <= "1110"; x_in <= "011000"; z_correct<="1111010000";
        when 903 => y_in <= "1111"; x_in <= "011000"; z_correct<="1111101000";
        when 904 => y_in <= "0000"; x_in <= "011000"; z_correct<="0000000000";
        when 905 => y_in <= "0001"; x_in <= "011000"; z_correct<="0000011000";
        when 906 => y_in <= "0010"; x_in <= "011000"; z_correct<="0000110000";
        when 907 => y_in <= "0011"; x_in <= "011000"; z_correct<="0001001000";
        when 908 => y_in <= "0100"; x_in <= "011000"; z_correct<="0001100000";
        when 909 => y_in <= "0101"; x_in <= "011000"; z_correct<="0001111000";
        when 910 => y_in <= "0110"; x_in <= "011000"; z_correct<="0010010000";
        when 911 => y_in <= "0111"; x_in <= "011000"; z_correct<="0010101000";
        when 912 => y_in <= "1000"; x_in <= "011001"; z_correct<="1100111000";
        when 913 => y_in <= "1001"; x_in <= "011001"; z_correct<="1101010001";
        when 914 => y_in <= "1010"; x_in <= "011001"; z_correct<="1101101010";
        when 915 => y_in <= "1011"; x_in <= "011001"; z_correct<="1110000011";
        when 916 => y_in <= "1100"; x_in <= "011001"; z_correct<="1110011100";
        when 917 => y_in <= "1101"; x_in <= "011001"; z_correct<="1110110101";
        when 918 => y_in <= "1110"; x_in <= "011001"; z_correct<="1111001110";
        when 919 => y_in <= "1111"; x_in <= "011001"; z_correct<="1111100111";
        when 920 => y_in <= "0000"; x_in <= "011001"; z_correct<="0000000000";
        when 921 => y_in <= "0001"; x_in <= "011001"; z_correct<="0000011001";
        when 922 => y_in <= "0010"; x_in <= "011001"; z_correct<="0000110010";
        when 923 => y_in <= "0011"; x_in <= "011001"; z_correct<="0001001011";
        when 924 => y_in <= "0100"; x_in <= "011001"; z_correct<="0001100100";
        when 925 => y_in <= "0101"; x_in <= "011001"; z_correct<="0001111101";
        when 926 => y_in <= "0110"; x_in <= "011001"; z_correct<="0010010110";
        when 927 => y_in <= "0111"; x_in <= "011001"; z_correct<="0010101111";
        when 928 => y_in <= "1000"; x_in <= "011010"; z_correct<="1100110000";
        when 929 => y_in <= "1001"; x_in <= "011010"; z_correct<="1101001010";
        when 930 => y_in <= "1010"; x_in <= "011010"; z_correct<="1101100100";
        when 931 => y_in <= "1011"; x_in <= "011010"; z_correct<="1101111110";
        when 932 => y_in <= "1100"; x_in <= "011010"; z_correct<="1110011000";
        when 933 => y_in <= "1101"; x_in <= "011010"; z_correct<="1110110010";
        when 934 => y_in <= "1110"; x_in <= "011010"; z_correct<="1111001100";
        when 935 => y_in <= "1111"; x_in <= "011010"; z_correct<="1111100110";
        when 936 => y_in <= "0000"; x_in <= "011010"; z_correct<="0000000000";
        when 937 => y_in <= "0001"; x_in <= "011010"; z_correct<="0000011010";
        when 938 => y_in <= "0010"; x_in <= "011010"; z_correct<="0000110100";
        when 939 => y_in <= "0011"; x_in <= "011010"; z_correct<="0001001110";
        when 940 => y_in <= "0100"; x_in <= "011010"; z_correct<="0001101000";
        when 941 => y_in <= "0101"; x_in <= "011010"; z_correct<="0010000010";
        when 942 => y_in <= "0110"; x_in <= "011010"; z_correct<="0010011100";
        when 943 => y_in <= "0111"; x_in <= "011010"; z_correct<="0010110110";
        when 944 => y_in <= "1000"; x_in <= "011011"; z_correct<="1100101000";
        when 945 => y_in <= "1001"; x_in <= "011011"; z_correct<="1101000011";
        when 946 => y_in <= "1010"; x_in <= "011011"; z_correct<="1101011110";
        when 947 => y_in <= "1011"; x_in <= "011011"; z_correct<="1101111001";
        when 948 => y_in <= "1100"; x_in <= "011011"; z_correct<="1110010100";
        when 949 => y_in <= "1101"; x_in <= "011011"; z_correct<="1110101111";
        when 950 => y_in <= "1110"; x_in <= "011011"; z_correct<="1111001010";
        when 951 => y_in <= "1111"; x_in <= "011011"; z_correct<="1111100101";
        when 952 => y_in <= "0000"; x_in <= "011011"; z_correct<="0000000000";
        when 953 => y_in <= "0001"; x_in <= "011011"; z_correct<="0000011011";
        when 954 => y_in <= "0010"; x_in <= "011011"; z_correct<="0000110110";
        when 955 => y_in <= "0011"; x_in <= "011011"; z_correct<="0001010001";
        when 956 => y_in <= "0100"; x_in <= "011011"; z_correct<="0001101100";
        when 957 => y_in <= "0101"; x_in <= "011011"; z_correct<="0010000111";
        when 958 => y_in <= "0110"; x_in <= "011011"; z_correct<="0010100010";
        when 959 => y_in <= "0111"; x_in <= "011011"; z_correct<="0010111101";
        when 960 => y_in <= "1000"; x_in <= "011100"; z_correct<="1100100000";
        when 961 => y_in <= "1001"; x_in <= "011100"; z_correct<="1100111100";
        when 962 => y_in <= "1010"; x_in <= "011100"; z_correct<="1101011000";
        when 963 => y_in <= "1011"; x_in <= "011100"; z_correct<="1101110100";
        when 964 => y_in <= "1100"; x_in <= "011100"; z_correct<="1110010000";
        when 965 => y_in <= "1101"; x_in <= "011100"; z_correct<="1110101100";
        when 966 => y_in <= "1110"; x_in <= "011100"; z_correct<="1111001000";
        when 967 => y_in <= "1111"; x_in <= "011100"; z_correct<="1111100100";
        when 968 => y_in <= "0000"; x_in <= "011100"; z_correct<="0000000000";
        when 969 => y_in <= "0001"; x_in <= "011100"; z_correct<="0000011100";
        when 970 => y_in <= "0010"; x_in <= "011100"; z_correct<="0000111000";
        when 971 => y_in <= "0011"; x_in <= "011100"; z_correct<="0001010100";
        when 972 => y_in <= "0100"; x_in <= "011100"; z_correct<="0001110000";
        when 973 => y_in <= "0101"; x_in <= "011100"; z_correct<="0010001100";
        when 974 => y_in <= "0110"; x_in <= "011100"; z_correct<="0010101000";
        when 975 => y_in <= "0111"; x_in <= "011100"; z_correct<="0011000100";
        when 976 => y_in <= "1000"; x_in <= "011101"; z_correct<="1100011000";
        when 977 => y_in <= "1001"; x_in <= "011101"; z_correct<="1100110101";
        when 978 => y_in <= "1010"; x_in <= "011101"; z_correct<="1101010010";
        when 979 => y_in <= "1011"; x_in <= "011101"; z_correct<="1101101111";
        when 980 => y_in <= "1100"; x_in <= "011101"; z_correct<="1110001100";
        when 981 => y_in <= "1101"; x_in <= "011101"; z_correct<="1110101001";
        when 982 => y_in <= "1110"; x_in <= "011101"; z_correct<="1111000110";
        when 983 => y_in <= "1111"; x_in <= "011101"; z_correct<="1111100011";
        when 984 => y_in <= "0000"; x_in <= "011101"; z_correct<="0000000000";
        when 985 => y_in <= "0001"; x_in <= "011101"; z_correct<="0000011101";
        when 986 => y_in <= "0010"; x_in <= "011101"; z_correct<="0000111010";
        when 987 => y_in <= "0011"; x_in <= "011101"; z_correct<="0001010111";
        when 988 => y_in <= "0100"; x_in <= "011101"; z_correct<="0001110100";
        when 989 => y_in <= "0101"; x_in <= "011101"; z_correct<="0010010001";
        when 990 => y_in <= "0110"; x_in <= "011101"; z_correct<="0010101110";
        when 991 => y_in <= "0111"; x_in <= "011101"; z_correct<="0011001011";
        when 992 => y_in <= "1000"; x_in <= "011110"; z_correct<="1100010000";
        when 993 => y_in <= "1001"; x_in <= "011110"; z_correct<="1100101110";
        when 994 => y_in <= "1010"; x_in <= "011110"; z_correct<="1101001100";
        when 995 => y_in <= "1011"; x_in <= "011110"; z_correct<="1101101010";
        when 996 => y_in <= "1100"; x_in <= "011110"; z_correct<="1110001000";
        when 997 => y_in <= "1101"; x_in <= "011110"; z_correct<="1110100110";
        when 998 => y_in <= "1110"; x_in <= "011110"; z_correct<="1111000100";
        when 999 => y_in <= "1111"; x_in <= "011110"; z_correct<="1111100010";
        when 1000 => y_in <= "0000"; x_in <= "011110"; z_correct<="0000000000";
        when 1001 => y_in <= "0001"; x_in <= "011110"; z_correct<="0000011110";
        when 1002 => y_in <= "0010"; x_in <= "011110"; z_correct<="0000111100";
        when 1003 => y_in <= "0011"; x_in <= "011110"; z_correct<="0001011010";
        when 1004 => y_in <= "0100"; x_in <= "011110"; z_correct<="0001111000";
        when 1005 => y_in <= "0101"; x_in <= "011110"; z_correct<="0010010110";
        when 1006 => y_in <= "0110"; x_in <= "011110"; z_correct<="0010110100";
        when 1007 => y_in <= "0111"; x_in <= "011110"; z_correct<="0011010010";
        when 1008 => y_in <= "1000"; x_in <= "011111"; z_correct<="1100001000";
        when 1009 => y_in <= "1001"; x_in <= "011111"; z_correct<="1100100111";
        when 1010 => y_in <= "1010"; x_in <= "011111"; z_correct<="1101000110";
        when 1011 => y_in <= "1011"; x_in <= "011111"; z_correct<="1101100101";
        when 1012 => y_in <= "1100"; x_in <= "011111"; z_correct<="1110000100";
        when 1013 => y_in <= "1101"; x_in <= "011111"; z_correct<="1110100011";
        when 1014 => y_in <= "1110"; x_in <= "011111"; z_correct<="1111000010";
        when 1015 => y_in <= "1111"; x_in <= "011111"; z_correct<="1111100001";
        when 1016 => y_in <= "0000"; x_in <= "011111"; z_correct<="0000000000";
        when 1017 => y_in <= "0001"; x_in <= "011111"; z_correct<="0000011111";
        when 1018 => y_in <= "0010"; x_in <= "011111"; z_correct<="0000111110";
        when 1019 => y_in <= "0011"; x_in <= "011111"; z_correct<="0001011101";
        when 1020 => y_in <= "0100"; x_in <= "011111"; z_correct<="0001111100";
        when 1021 => y_in <= "0101"; x_in <= "011111"; z_correct<="0010011011";
        when 1022 => y_in <= "0110"; x_in <= "011111"; z_correct<="0010111010";
        when 1023 => y_in <= "0111"; x_in <= "011111"; z_correct<="0011011001";

        when 1024 =>   Testing <= False;
        when others => null;
     end case;
	 if (z_out = z_correct) then diff <= '0'; else diff <= '1'; end if;
     count:= count + 1;
   end process Test_Proc;
end booth2_tbnm;
