

library IEEE;
use IEEE.std_logic_1164.all;

entity booth2_tbn4 IS

end booth2_tbn4;

-- Test Booth Multiplier with N=M=4

architecture booth2_tbn4 of booth2_tbn4 is
	component Booth2Multiplier
  	generic(N : integer := 4; 
            M : integer := 4   
       );
	port (
	x : in  std_logic_vector(N-1 downto 0); 	-- x is the multiplicand
	y : in  std_logic_vector(M-1 downto 0);		-- y is the multiplier
	z : out	std_logic_vector(N+M-1 downto 0)	-- z is the result of the multiplication
		);
	end component; 
	
   constant MckPer  :  time     := 200 ns; 
	   
   signal   clk  : std_logic := '0';
   signal   x_in   	: std_logic_VECTOR (3 downto 0):="0000";
   signal   y_in    : std_logic_VECTOR (3 downto 0):="0000";	
   signal   z_out   : std_logic_VECTOR (7 downto 0):="00000000";
   signal clk_cycle : integer;
   signal Testing: boolean := True;	
   signal z_correct   : std_logic_VECTOR (7 downto 0):="00000000";
   signal 	diff		: std_logic := '0';
begin 			 
	I: Booth2Multiplier generic map(N=>4, M=>4)
		port map(x=>x_in,y=>y_in, z=>z_out);
				
		clk <= not clk after MckPer/2 when Testing else '0';


   Test_Proc: process(clk)
   variable count: INTEGER:= 0;
   
   begin
     clk_cycle <= (count+1)/2;

     case clk_cycle is
        when 0 => y_in <= "1000"; x_in <= "1000"; z_correct<="01000000";
        when 1 => y_in <= "1000"; x_in <= "1001"; z_correct<="00111000";
        when 2 => y_in <= "1000"; x_in <= "1010"; z_correct<="00110000";
        when 3 => y_in <= "1000"; x_in <= "1011"; z_correct<="00101000";
        when 4 => y_in <= "1000"; x_in <= "1100"; z_correct<="00100000";
        when 5 => y_in <= "1000"; x_in <= "1101"; z_correct<="00011000";
        when 6 => y_in <= "1000"; x_in <= "1110"; z_correct<="00010000";
        when 7 => y_in <= "1000"; x_in <= "1111"; z_correct<="00001000";
        when 8 => y_in <= "1000"; x_in <= "0000"; z_correct<="00000000";
        when 9 => y_in <= "1000"; x_in <= "0001"; z_correct<="11111000";
        when 10 => y_in <= "1000"; x_in <= "0010"; z_correct<="11110000";
        when 11 => y_in <= "1000"; x_in <= "0011"; z_correct<="11101000";
        when 12 => y_in <= "1000"; x_in <= "0100"; z_correct<="11100000";
        when 13 => y_in <= "1000"; x_in <= "0101"; z_correct<="11011000";
        when 14 => y_in <= "1000"; x_in <= "0110"; z_correct<="11010000";
        when 15 => y_in <= "1000"; x_in <= "0111"; z_correct<="11001000";
        when 16 => y_in <= "1001"; x_in <= "1000"; z_correct<="00111000";
        when 17 => y_in <= "1001"; x_in <= "1001"; z_correct<="00110001";
        when 18 => y_in <= "1001"; x_in <= "1010"; z_correct<="00101010";
        when 19 => y_in <= "1001"; x_in <= "1011"; z_correct<="00100011";
        when 20 => y_in <= "1001"; x_in <= "1100"; z_correct<="00011100";
        when 21 => y_in <= "1001"; x_in <= "1101"; z_correct<="00010101";
        when 22 => y_in <= "1001"; x_in <= "1110"; z_correct<="00001110";
        when 23 => y_in <= "1001"; x_in <= "1111"; z_correct<="00000111";
        when 24 => y_in <= "1001"; x_in <= "0000"; z_correct<="00000000";
        when 25 => y_in <= "1001"; x_in <= "0001"; z_correct<="11111001";
        when 26 => y_in <= "1001"; x_in <= "0010"; z_correct<="11110010";
        when 27 => y_in <= "1001"; x_in <= "0011"; z_correct<="11101011";
        when 28 => y_in <= "1001"; x_in <= "0100"; z_correct<="11100100";
        when 29 => y_in <= "1001"; x_in <= "0101"; z_correct<="11011101";
        when 30 => y_in <= "1001"; x_in <= "0110"; z_correct<="11010110";
        when 31 => y_in <= "1001"; x_in <= "0111"; z_correct<="11001111";
        when 32 => y_in <= "1010"; x_in <= "1000"; z_correct<="00110000";
        when 33 => y_in <= "1010"; x_in <= "1001"; z_correct<="00101010";
        when 34 => y_in <= "1010"; x_in <= "1010"; z_correct<="00100100";
        when 35 => y_in <= "1010"; x_in <= "1011"; z_correct<="00011110";
        when 36 => y_in <= "1010"; x_in <= "1100"; z_correct<="00011000";
        when 37 => y_in <= "1010"; x_in <= "1101"; z_correct<="00010010";
        when 38 => y_in <= "1010"; x_in <= "1110"; z_correct<="00001100";
        when 39 => y_in <= "1010"; x_in <= "1111"; z_correct<="00000110";
        when 40 => y_in <= "1010"; x_in <= "0000"; z_correct<="00000000";
        when 41 => y_in <= "1010"; x_in <= "0001"; z_correct<="11111010";
        when 42 => y_in <= "1010"; x_in <= "0010"; z_correct<="11110100";
        when 43 => y_in <= "1010"; x_in <= "0011"; z_correct<="11101110";
        when 44 => y_in <= "1010"; x_in <= "0100"; z_correct<="11101000";
        when 45 => y_in <= "1010"; x_in <= "0101"; z_correct<="11100010";
        when 46 => y_in <= "1010"; x_in <= "0110"; z_correct<="11011100";
        when 47 => y_in <= "1010"; x_in <= "0111"; z_correct<="11010110";
        when 48 => y_in <= "1011"; x_in <= "1000"; z_correct<="00101000";
        when 49 => y_in <= "1011"; x_in <= "1001"; z_correct<="00100011";
        when 50 => y_in <= "1011"; x_in <= "1010"; z_correct<="00011110";
        when 51 => y_in <= "1011"; x_in <= "1011"; z_correct<="00011001";
        when 52 => y_in <= "1011"; x_in <= "1100"; z_correct<="00010100";
        when 53 => y_in <= "1011"; x_in <= "1101"; z_correct<="00001111";
        when 54 => y_in <= "1011"; x_in <= "1110"; z_correct<="00001010";
        when 55 => y_in <= "1011"; x_in <= "1111"; z_correct<="00000101";
        when 56 => y_in <= "1011"; x_in <= "0000"; z_correct<="00000000";
        when 57 => y_in <= "1011"; x_in <= "0001"; z_correct<="11111011";
        when 58 => y_in <= "1011"; x_in <= "0010"; z_correct<="11110110";
        when 59 => y_in <= "1011"; x_in <= "0011"; z_correct<="11110001";
        when 60 => y_in <= "1011"; x_in <= "0100"; z_correct<="11101100";
        when 61 => y_in <= "1011"; x_in <= "0101"; z_correct<="11100111";
        when 62 => y_in <= "1011"; x_in <= "0110"; z_correct<="11100010";
        when 63 => y_in <= "1011"; x_in <= "0111"; z_correct<="11011101";
        when 64 => y_in <= "1100"; x_in <= "1000"; z_correct<="00100000";
        when 65 => y_in <= "1100"; x_in <= "1001"; z_correct<="00011100";
        when 66 => y_in <= "1100"; x_in <= "1010"; z_correct<="00011000";
        when 67 => y_in <= "1100"; x_in <= "1011"; z_correct<="00010100";
        when 68 => y_in <= "1100"; x_in <= "1100"; z_correct<="00010000";
        when 69 => y_in <= "1100"; x_in <= "1101"; z_correct<="00001100";
        when 70 => y_in <= "1100"; x_in <= "1110"; z_correct<="00001000";
        when 71 => y_in <= "1100"; x_in <= "1111"; z_correct<="00000100";
        when 72 => y_in <= "1100"; x_in <= "0000"; z_correct<="00000000";
        when 73 => y_in <= "1100"; x_in <= "0001"; z_correct<="11111100";
        when 74 => y_in <= "1100"; x_in <= "0010"; z_correct<="11111000";
        when 75 => y_in <= "1100"; x_in <= "0011"; z_correct<="11110100";
        when 76 => y_in <= "1100"; x_in <= "0100"; z_correct<="11110000";
        when 77 => y_in <= "1100"; x_in <= "0101"; z_correct<="11101100";
        when 78 => y_in <= "1100"; x_in <= "0110"; z_correct<="11101000";
        when 79 => y_in <= "1100"; x_in <= "0111"; z_correct<="11100100";
        when 80 => y_in <= "1101"; x_in <= "1000"; z_correct<="00011000";
        when 81 => y_in <= "1101"; x_in <= "1001"; z_correct<="00010101";
        when 82 => y_in <= "1101"; x_in <= "1010"; z_correct<="00010010";
        when 83 => y_in <= "1101"; x_in <= "1011"; z_correct<="00001111";
        when 84 => y_in <= "1101"; x_in <= "1100"; z_correct<="00001100";
        when 85 => y_in <= "1101"; x_in <= "1101"; z_correct<="00001001";
        when 86 => y_in <= "1101"; x_in <= "1110"; z_correct<="00000110";
        when 87 => y_in <= "1101"; x_in <= "1111"; z_correct<="00000011";
        when 88 => y_in <= "1101"; x_in <= "0000"; z_correct<="00000000";
        when 89 => y_in <= "1101"; x_in <= "0001"; z_correct<="11111101";
        when 90 => y_in <= "1101"; x_in <= "0010"; z_correct<="11111010";
        when 91 => y_in <= "1101"; x_in <= "0011"; z_correct<="11110111";
        when 92 => y_in <= "1101"; x_in <= "0100"; z_correct<="11110100";
        when 93 => y_in <= "1101"; x_in <= "0101"; z_correct<="11110001";
        when 94 => y_in <= "1101"; x_in <= "0110"; z_correct<="11101110";
        when 95 => y_in <= "1101"; x_in <= "0111"; z_correct<="11101011";
        when 96 => y_in <= "1110"; x_in <= "1000"; z_correct<="00010000";
        when 97 => y_in <= "1110"; x_in <= "1001"; z_correct<="00001110";
        when 98 => y_in <= "1110"; x_in <= "1010"; z_correct<="00001100";
        when 99 => y_in <= "1110"; x_in <= "1011"; z_correct<="00001010";
        when 100 => y_in <= "1110"; x_in <= "1100"; z_correct<="00001000";
        when 101 => y_in <= "1110"; x_in <= "1101"; z_correct<="00000110";
        when 102 => y_in <= "1110"; x_in <= "1110"; z_correct<="00000100";
        when 103 => y_in <= "1110"; x_in <= "1111"; z_correct<="00000010";
        when 104 => y_in <= "1110"; x_in <= "0000"; z_correct<="00000000";
        when 105 => y_in <= "1110"; x_in <= "0001"; z_correct<="11111110";
        when 106 => y_in <= "1110"; x_in <= "0010"; z_correct<="11111100";
        when 107 => y_in <= "1110"; x_in <= "0011"; z_correct<="11111010";
        when 108 => y_in <= "1110"; x_in <= "0100"; z_correct<="11111000";
        when 109 => y_in <= "1110"; x_in <= "0101"; z_correct<="11110110";
        when 110 => y_in <= "1110"; x_in <= "0110"; z_correct<="11110100";
        when 111 => y_in <= "1110"; x_in <= "0111"; z_correct<="11110010";
        when 112 => y_in <= "1111"; x_in <= "1000"; z_correct<="00001000";
        when 113 => y_in <= "1111"; x_in <= "1001"; z_correct<="00000111";
        when 114 => y_in <= "1111"; x_in <= "1010"; z_correct<="00000110";
        when 115 => y_in <= "1111"; x_in <= "1011"; z_correct<="00000101";
        when 116 => y_in <= "1111"; x_in <= "1100"; z_correct<="00000100";
        when 117 => y_in <= "1111"; x_in <= "1101"; z_correct<="00000011";
        when 118 => y_in <= "1111"; x_in <= "1110"; z_correct<="00000010";
        when 119 => y_in <= "1111"; x_in <= "1111"; z_correct<="00000001";
        when 120 => y_in <= "1111"; x_in <= "0000"; z_correct<="00000000";
        when 121 => y_in <= "1111"; x_in <= "0001"; z_correct<="11111111";
        when 122 => y_in <= "1111"; x_in <= "0010"; z_correct<="11111110";
        when 123 => y_in <= "1111"; x_in <= "0011"; z_correct<="11111101";
        when 124 => y_in <= "1111"; x_in <= "0100"; z_correct<="11111100";
        when 125 => y_in <= "1111"; x_in <= "0101"; z_correct<="11111011";
        when 126 => y_in <= "1111"; x_in <= "0110"; z_correct<="11111010";
        when 127 => y_in <= "1111"; x_in <= "0111"; z_correct<="11111001";
        when 128 => y_in <= "0000"; x_in <= "1000"; z_correct<="00000000";
        when 129 => y_in <= "0000"; x_in <= "1001"; z_correct<="00000000";
        when 130 => y_in <= "0000"; x_in <= "1010"; z_correct<="00000000";
        when 131 => y_in <= "0000"; x_in <= "1011"; z_correct<="00000000";
        when 132 => y_in <= "0000"; x_in <= "1100"; z_correct<="00000000";
        when 133 => y_in <= "0000"; x_in <= "1101"; z_correct<="00000000";
        when 134 => y_in <= "0000"; x_in <= "1110"; z_correct<="00000000";
        when 135 => y_in <= "0000"; x_in <= "1111"; z_correct<="00000000";
        when 136 => y_in <= "0000"; x_in <= "0000"; z_correct<="00000000";
        when 137 => y_in <= "0000"; x_in <= "0001"; z_correct<="00000000";
        when 138 => y_in <= "0000"; x_in <= "0010"; z_correct<="00000000";
        when 139 => y_in <= "0000"; x_in <= "0011"; z_correct<="00000000";
        when 140 => y_in <= "0000"; x_in <= "0100"; z_correct<="00000000";
        when 141 => y_in <= "0000"; x_in <= "0101"; z_correct<="00000000";
        when 142 => y_in <= "0000"; x_in <= "0110"; z_correct<="00000000";
        when 143 => y_in <= "0000"; x_in <= "0111"; z_correct<="00000000";
        when 144 => y_in <= "0001"; x_in <= "1000"; z_correct<="11111000";
        when 145 => y_in <= "0001"; x_in <= "1001"; z_correct<="11111001";
        when 146 => y_in <= "0001"; x_in <= "1010"; z_correct<="11111010";
        when 147 => y_in <= "0001"; x_in <= "1011"; z_correct<="11111011";
        when 148 => y_in <= "0001"; x_in <= "1100"; z_correct<="11111100";
        when 149 => y_in <= "0001"; x_in <= "1101"; z_correct<="11111101";
        when 150 => y_in <= "0001"; x_in <= "1110"; z_correct<="11111110";
        when 151 => y_in <= "0001"; x_in <= "1111"; z_correct<="11111111";
        when 152 => y_in <= "0001"; x_in <= "0000"; z_correct<="00000000";
        when 153 => y_in <= "0001"; x_in <= "0001"; z_correct<="00000001";
        when 154 => y_in <= "0001"; x_in <= "0010"; z_correct<="00000010";
        when 155 => y_in <= "0001"; x_in <= "0011"; z_correct<="00000011";
        when 156 => y_in <= "0001"; x_in <= "0100"; z_correct<="00000100";
        when 157 => y_in <= "0001"; x_in <= "0101"; z_correct<="00000101";
        when 158 => y_in <= "0001"; x_in <= "0110"; z_correct<="00000110";
        when 159 => y_in <= "0001"; x_in <= "0111"; z_correct<="00000111";
        when 160 => y_in <= "0010"; x_in <= "1000"; z_correct<="11110000";
        when 161 => y_in <= "0010"; x_in <= "1001"; z_correct<="11110010";
        when 162 => y_in <= "0010"; x_in <= "1010"; z_correct<="11110100";
        when 163 => y_in <= "0010"; x_in <= "1011"; z_correct<="11110110";
        when 164 => y_in <= "0010"; x_in <= "1100"; z_correct<="11111000";
        when 165 => y_in <= "0010"; x_in <= "1101"; z_correct<="11111010";
        when 166 => y_in <= "0010"; x_in <= "1110"; z_correct<="11111100";
        when 167 => y_in <= "0010"; x_in <= "1111"; z_correct<="11111110";
        when 168 => y_in <= "0010"; x_in <= "0000"; z_correct<="00000000";
        when 169 => y_in <= "0010"; x_in <= "0001"; z_correct<="00000010";
        when 170 => y_in <= "0010"; x_in <= "0010"; z_correct<="00000100";
        when 171 => y_in <= "0010"; x_in <= "0011"; z_correct<="00000110";
        when 172 => y_in <= "0010"; x_in <= "0100"; z_correct<="00001000";
        when 173 => y_in <= "0010"; x_in <= "0101"; z_correct<="00001010";
        when 174 => y_in <= "0010"; x_in <= "0110"; z_correct<="00001100";
        when 175 => y_in <= "0010"; x_in <= "0111"; z_correct<="00001110";
        when 176 => y_in <= "0011"; x_in <= "1000"; z_correct<="11101000";
        when 177 => y_in <= "0011"; x_in <= "1001"; z_correct<="11101011";
        when 178 => y_in <= "0011"; x_in <= "1010"; z_correct<="11101110";
        when 179 => y_in <= "0011"; x_in <= "1011"; z_correct<="11110001";
        when 180 => y_in <= "0011"; x_in <= "1100"; z_correct<="11110100";
        when 181 => y_in <= "0011"; x_in <= "1101"; z_correct<="11110111";
        when 182 => y_in <= "0011"; x_in <= "1110"; z_correct<="11111010";
        when 183 => y_in <= "0011"; x_in <= "1111"; z_correct<="11111101";
        when 184 => y_in <= "0011"; x_in <= "0000"; z_correct<="00000000";
        when 185 => y_in <= "0011"; x_in <= "0001"; z_correct<="00000011";
        when 186 => y_in <= "0011"; x_in <= "0010"; z_correct<="00000110";
        when 187 => y_in <= "0011"; x_in <= "0011"; z_correct<="00001001";
        when 188 => y_in <= "0011"; x_in <= "0100"; z_correct<="00001100";
        when 189 => y_in <= "0011"; x_in <= "0101"; z_correct<="00001111";
        when 190 => y_in <= "0011"; x_in <= "0110"; z_correct<="00010010";
        when 191 => y_in <= "0011"; x_in <= "0111"; z_correct<="00010101";
        when 192 => y_in <= "0100"; x_in <= "1000"; z_correct<="11100000";
        when 193 => y_in <= "0100"; x_in <= "1001"; z_correct<="11100100";
        when 194 => y_in <= "0100"; x_in <= "1010"; z_correct<="11101000";
        when 195 => y_in <= "0100"; x_in <= "1011"; z_correct<="11101100";
        when 196 => y_in <= "0100"; x_in <= "1100"; z_correct<="11110000";
        when 197 => y_in <= "0100"; x_in <= "1101"; z_correct<="11110100";
        when 198 => y_in <= "0100"; x_in <= "1110"; z_correct<="11111000";
        when 199 => y_in <= "0100"; x_in <= "1111"; z_correct<="11111100";
        when 200 => y_in <= "0100"; x_in <= "0000"; z_correct<="00000000";
        when 201 => y_in <= "0100"; x_in <= "0001"; z_correct<="00000100";
        when 202 => y_in <= "0100"; x_in <= "0010"; z_correct<="00001000";
        when 203 => y_in <= "0100"; x_in <= "0011"; z_correct<="00001100";
        when 204 => y_in <= "0100"; x_in <= "0100"; z_correct<="00010000";
        when 205 => y_in <= "0100"; x_in <= "0101"; z_correct<="00010100";
        when 206 => y_in <= "0100"; x_in <= "0110"; z_correct<="00011000";
        when 207 => y_in <= "0100"; x_in <= "0111"; z_correct<="00011100";
        when 208 => y_in <= "0101"; x_in <= "1000"; z_correct<="11011000";
        when 209 => y_in <= "0101"; x_in <= "1001"; z_correct<="11011101";
        when 210 => y_in <= "0101"; x_in <= "1010"; z_correct<="11100010";
        when 211 => y_in <= "0101"; x_in <= "1011"; z_correct<="11100111";
        when 212 => y_in <= "0101"; x_in <= "1100"; z_correct<="11101100";
        when 213 => y_in <= "0101"; x_in <= "1101"; z_correct<="11110001";
        when 214 => y_in <= "0101"; x_in <= "1110"; z_correct<="11110110";
        when 215 => y_in <= "0101"; x_in <= "1111"; z_correct<="11111011";
        when 216 => y_in <= "0101"; x_in <= "0000"; z_correct<="00000000";
        when 217 => y_in <= "0101"; x_in <= "0001"; z_correct<="00000101";
        when 218 => y_in <= "0101"; x_in <= "0010"; z_correct<="00001010";
        when 219 => y_in <= "0101"; x_in <= "0011"; z_correct<="00001111";
        when 220 => y_in <= "0101"; x_in <= "0100"; z_correct<="00010100";
        when 221 => y_in <= "0101"; x_in <= "0101"; z_correct<="00011001";
        when 222 => y_in <= "0101"; x_in <= "0110"; z_correct<="00011110";
        when 223 => y_in <= "0101"; x_in <= "0111"; z_correct<="00100011";
        when 224 => y_in <= "0110"; x_in <= "1000"; z_correct<="11010000";
        when 225 => y_in <= "0110"; x_in <= "1001"; z_correct<="11010110";
        when 226 => y_in <= "0110"; x_in <= "1010"; z_correct<="11011100";
        when 227 => y_in <= "0110"; x_in <= "1011"; z_correct<="11100010";
        when 228 => y_in <= "0110"; x_in <= "1100"; z_correct<="11101000";
        when 229 => y_in <= "0110"; x_in <= "1101"; z_correct<="11101110";
        when 230 => y_in <= "0110"; x_in <= "1110"; z_correct<="11110100";
        when 231 => y_in <= "0110"; x_in <= "1111"; z_correct<="11111010";
        when 232 => y_in <= "0110"; x_in <= "0000"; z_correct<="00000000";
        when 233 => y_in <= "0110"; x_in <= "0001"; z_correct<="00000110";
        when 234 => y_in <= "0110"; x_in <= "0010"; z_correct<="00001100";
        when 235 => y_in <= "0110"; x_in <= "0011"; z_correct<="00010010";
        when 236 => y_in <= "0110"; x_in <= "0100"; z_correct<="00011000";
        when 237 => y_in <= "0110"; x_in <= "0101"; z_correct<="00011110";
        when 238 => y_in <= "0110"; x_in <= "0110"; z_correct<="00100100";
        when 239 => y_in <= "0110"; x_in <= "0111"; z_correct<="00101010";
        when 240 => y_in <= "0111"; x_in <= "1000"; z_correct<="11001000";
        when 241 => y_in <= "0111"; x_in <= "1001"; z_correct<="11001111";
        when 242 => y_in <= "0111"; x_in <= "1010"; z_correct<="11010110";
        when 243 => y_in <= "0111"; x_in <= "1011"; z_correct<="11011101";
        when 244 => y_in <= "0111"; x_in <= "1100"; z_correct<="11100100";
        when 245 => y_in <= "0111"; x_in <= "1101"; z_correct<="11101011";
        when 246 => y_in <= "0111"; x_in <= "1110"; z_correct<="11110010";
        when 247 => y_in <= "0111"; x_in <= "1111"; z_correct<="11111001";
        when 248 => y_in <= "0111"; x_in <= "0000"; z_correct<="00000000";
        when 249 => y_in <= "0111"; x_in <= "0001"; z_correct<="00000111";
        when 250 => y_in <= "0111"; x_in <= "0010"; z_correct<="00001110";
        when 251 => y_in <= "0111"; x_in <= "0011"; z_correct<="00010101";
        when 252 => y_in <= "0111"; x_in <= "0100"; z_correct<="00011100";
        when 253 => y_in <= "0111"; x_in <= "0101"; z_correct<="00100011";
        when 254 => y_in <= "0111"; x_in <= "0110"; z_correct<="00101010";
        when 255 => y_in <= "0111"; x_in <= "0111"; z_correct<="00110001";

        when 256 =>   Testing <= False;
        when others => null;
     end case;
	 if (z_out = z_correct) then diff <= '0'; else diff <= '1'; end if;
     count:= count + 1;
   end process Test_Proc;
end booth2_tbn4;
